-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bbd",
     9 => x"e0080b0b",
    10 => x"0bbde408",
    11 => x"0b0b0bbd",
    12 => x"e8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bde80c0b",
    16 => x"0b0bbde4",
    17 => x"0c0b0b0b",
    18 => x"bde00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb28c",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bde07080",
    57 => x"c890278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188e304",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbdf00c",
    65 => x"9f0bbdf4",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bdf408ff",
    69 => x"05bdf40c",
    70 => x"bdf40880",
    71 => x"25eb38bd",
    72 => x"f008ff05",
    73 => x"bdf00cbd",
    74 => x"f0088025",
    75 => x"d738800b",
    76 => x"bdf40c80",
    77 => x"0bbdf00c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bbdf008",
    97 => x"258f3882",
    98 => x"bd2dbdf0",
    99 => x"08ff05bd",
   100 => x"f00c82ff",
   101 => x"04bdf008",
   102 => x"bdf40853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"bdf008a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134bdf4",
   111 => x"088105bd",
   112 => x"f40cbdf4",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bbdf40c",
   116 => x"bdf00881",
   117 => x"05bdf00c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134bd",
   122 => x"f4088105",
   123 => x"bdf40cbd",
   124 => x"f408a02e",
   125 => x"0981068e",
   126 => x"38800bbd",
   127 => x"f40cbdf0",
   128 => x"088105bd",
   129 => x"f00c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bbdf8",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bbdf80c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872bd",
   169 => x"f8088407",
   170 => x"bdf80c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb8e8",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"bdf80852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"bde00c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dec51",
   218 => x"92710c86",
   219 => x"a42d8271",
   220 => x"0c028405",
   221 => x"0d0402d0",
   222 => x"050d7d54",
   223 => x"805ba40b",
   224 => x"ec0c7352",
   225 => x"bdfc51a9",
   226 => x"ac2dbde0",
   227 => x"087b2e81",
   228 => x"ab38be80",
   229 => x"0870f80c",
   230 => x"891580f5",
   231 => x"2d8a1680",
   232 => x"f52d7182",
   233 => x"80290588",
   234 => x"1780f52d",
   235 => x"70848080",
   236 => x"2912f40c",
   237 => x"7eff155c",
   238 => x"5e575556",
   239 => x"58767b2e",
   240 => x"8b38811a",
   241 => x"77812a58",
   242 => x"5a76f738",
   243 => x"f71a5a81",
   244 => x"5b807825",
   245 => x"80e63879",
   246 => x"52765184",
   247 => x"8b2dbec8",
   248 => x"52bdfc51",
   249 => x"abeb2dbd",
   250 => x"e008802e",
   251 => x"b838bec8",
   252 => x"5c83fc59",
   253 => x"7b708405",
   254 => x"5d087081",
   255 => x"ff067188",
   256 => x"2a7081ff",
   257 => x"0673902a",
   258 => x"7081ff06",
   259 => x"75982ae8",
   260 => x"0ce80c58",
   261 => x"e80c57e8",
   262 => x"0cfc1a5a",
   263 => x"53788025",
   264 => x"d33888ac",
   265 => x"04bde008",
   266 => x"5b848058",
   267 => x"bdfc51ab",
   268 => x"bd2dfc80",
   269 => x"18811858",
   270 => x"5887d104",
   271 => x"86b72d84",
   272 => x"0bec0c7a",
   273 => x"802e8d38",
   274 => x"b8ec5191",
   275 => x"d22d8fd5",
   276 => x"2d88da04",
   277 => x"bbb05191",
   278 => x"d22d7abd",
   279 => x"e00c02b0",
   280 => x"050d0402",
   281 => x"d4050d80",
   282 => x"55840bec",
   283 => x"0c8fb62d",
   284 => x"8ca02d81",
   285 => x"f82da0a1",
   286 => x"2dbde008",
   287 => x"752e838b",
   288 => x"388c0bec",
   289 => x"0cb7a852",
   290 => x"bdfc51a9",
   291 => x"ac2dbde0",
   292 => x"08752e81",
   293 => x"8338be80",
   294 => x"0875ff12",
   295 => x"595b5876",
   296 => x"752e8b38",
   297 => x"811a7781",
   298 => x"2a585a76",
   299 => x"f738f71a",
   300 => x"5a807825",
   301 => x"80e23879",
   302 => x"52765184",
   303 => x"8b2dbec8",
   304 => x"52bdfc51",
   305 => x"abeb2dbd",
   306 => x"e008802e",
   307 => x"b838bec8",
   308 => x"5b83fc59",
   309 => x"7a708405",
   310 => x"5c087081",
   311 => x"ff067188",
   312 => x"2a7081ff",
   313 => x"0673902a",
   314 => x"7081ff06",
   315 => x"75982ae8",
   316 => x"0ce80c58",
   317 => x"e80c57e8",
   318 => x"0cfc1a5a",
   319 => x"53788025",
   320 => x"d3388a88",
   321 => x"04848058",
   322 => x"bdfc51ab",
   323 => x"bd2dfc80",
   324 => x"18811858",
   325 => x"5889b104",
   326 => x"be8008f8",
   327 => x"0c86b72d",
   328 => x"840bec0c",
   329 => x"86f651b2",
   330 => x"852db8ec",
   331 => x"5191d22d",
   332 => x"8fd52d8c",
   333 => x"ac2d91e2",
   334 => x"2db9800b",
   335 => x"80f52d70",
   336 => x"862b80c0",
   337 => x"06b98c0b",
   338 => x"80f52d70",
   339 => x"872b8180",
   340 => x"06b9980b",
   341 => x"80f52d70",
   342 => x"852ba006",
   343 => x"74730707",
   344 => x"b9a40b80",
   345 => x"f52d708c",
   346 => x"2b80e080",
   347 => x"06b9b00b",
   348 => x"80f52d70",
   349 => x"842b9006",
   350 => x"74730707",
   351 => x"b9bc0b80",
   352 => x"f52d7091",
   353 => x"2b988080",
   354 => x"06b9c80b",
   355 => x"80f52d70",
   356 => x"8a2b9880",
   357 => x"06747307",
   358 => x"07b9d40b",
   359 => x"80f52d70",
   360 => x"902b8480",
   361 => x"8006b9e0",
   362 => x"0b80f52d",
   363 => x"708e2b83",
   364 => x"80800674",
   365 => x"730707b9",
   366 => x"ec0b80f5",
   367 => x"2d70932b",
   368 => x"a0808006",
   369 => x"b9f80b80",
   370 => x"f52d7094",
   371 => x"2b90800a",
   372 => x"06747307",
   373 => x"07ba840b",
   374 => x"80f52d70",
   375 => x"882b8680",
   376 => x"067207fc",
   377 => x"0c535454",
   378 => x"54545454",
   379 => x"54545454",
   380 => x"54545454",
   381 => x"54565452",
   382 => x"57585653",
   383 => x"8653bde0",
   384 => x"08833884",
   385 => x"5372ec0c",
   386 => x"8ab30480",
   387 => x"0bbde00c",
   388 => x"02ac050d",
   389 => x"0471980c",
   390 => x"04ffb008",
   391 => x"bde00c04",
   392 => x"810bffb0",
   393 => x"0c04800b",
   394 => x"ffb00c04",
   395 => x"02f4050d",
   396 => x"8dae04bd",
   397 => x"e00881f0",
   398 => x"2e098106",
   399 => x"8938810b",
   400 => x"bc940c8d",
   401 => x"ae04bde0",
   402 => x"0881e02e",
   403 => x"09810689",
   404 => x"38810bbc",
   405 => x"980c8dae",
   406 => x"04bde008",
   407 => x"52bc9808",
   408 => x"802e8838",
   409 => x"bde00881",
   410 => x"80055271",
   411 => x"842c728f",
   412 => x"065353bc",
   413 => x"9408802e",
   414 => x"99387284",
   415 => x"29bbd405",
   416 => x"72138171",
   417 => x"2b700973",
   418 => x"0806730c",
   419 => x"5153538d",
   420 => x"a4047284",
   421 => x"29bbd405",
   422 => x"72138371",
   423 => x"2b720807",
   424 => x"720c5353",
   425 => x"800bbc98",
   426 => x"0c800bbc",
   427 => x"940cbe88",
   428 => x"518eaf2d",
   429 => x"bde008ff",
   430 => x"24fef838",
   431 => x"800bbde0",
   432 => x"0c028c05",
   433 => x"0d0402f8",
   434 => x"050dbbd4",
   435 => x"528f5180",
   436 => x"72708405",
   437 => x"540cff11",
   438 => x"51708025",
   439 => x"f2380288",
   440 => x"050d0402",
   441 => x"f0050d75",
   442 => x"518ca62d",
   443 => x"70822cfc",
   444 => x"06bbd411",
   445 => x"72109e06",
   446 => x"71087072",
   447 => x"2a708306",
   448 => x"82742b70",
   449 => x"09740676",
   450 => x"0c545156",
   451 => x"57535153",
   452 => x"8ca02d71",
   453 => x"bde00c02",
   454 => x"90050d04",
   455 => x"02fc050d",
   456 => x"72518071",
   457 => x"0c800b84",
   458 => x"120c0284",
   459 => x"050d0402",
   460 => x"f0050d75",
   461 => x"70088412",
   462 => x"08535353",
   463 => x"ff547171",
   464 => x"2ea8388c",
   465 => x"a62d8413",
   466 => x"08708429",
   467 => x"14881170",
   468 => x"087081ff",
   469 => x"06841808",
   470 => x"81118706",
   471 => x"841a0c53",
   472 => x"51555151",
   473 => x"518ca02d",
   474 => x"715473bd",
   475 => x"e00c0290",
   476 => x"050d0402",
   477 => x"f8050d8c",
   478 => x"a62de008",
   479 => x"708b2a70",
   480 => x"81065152",
   481 => x"5270802e",
   482 => x"9d38be88",
   483 => x"08708429",
   484 => x"be900573",
   485 => x"81ff0671",
   486 => x"0c5151be",
   487 => x"88088111",
   488 => x"8706be88",
   489 => x"0c51800b",
   490 => x"beb00c8c",
   491 => x"992d8ca0",
   492 => x"2d028805",
   493 => x"0d0402fc",
   494 => x"050dbe88",
   495 => x"518e9c2d",
   496 => x"8dc62d8e",
   497 => x"f3518c95",
   498 => x"2d028405",
   499 => x"0d04beb4",
   500 => x"08bde00c",
   501 => x"0402fc05",
   502 => x"0d8fdf04",
   503 => x"8cac2d80",
   504 => x"f6518de3",
   505 => x"2dbde008",
   506 => x"f33880da",
   507 => x"518de32d",
   508 => x"bde008e8",
   509 => x"38bde008",
   510 => x"bca00cbd",
   511 => x"e0085184",
   512 => x"f02d0284",
   513 => x"050d0402",
   514 => x"ec050d76",
   515 => x"54805287",
   516 => x"0b881580",
   517 => x"f52d5653",
   518 => x"74722483",
   519 => x"38a05372",
   520 => x"5182f92d",
   521 => x"81128b15",
   522 => x"80f52d54",
   523 => x"52727225",
   524 => x"de380294",
   525 => x"050d0402",
   526 => x"f0050dbe",
   527 => x"b4085481",
   528 => x"f82d800b",
   529 => x"beb80c73",
   530 => x"08802e81",
   531 => x"8038820b",
   532 => x"bdf40cbe",
   533 => x"b8088f06",
   534 => x"bdf00c73",
   535 => x"08527183",
   536 => x"2e963871",
   537 => x"83268938",
   538 => x"71812eaf",
   539 => x"3891b804",
   540 => x"71852e9f",
   541 => x"3891b804",
   542 => x"881480f5",
   543 => x"2d841508",
   544 => x"b7b45354",
   545 => x"5285fe2d",
   546 => x"71842913",
   547 => x"70085252",
   548 => x"91bc0473",
   549 => x"5190872d",
   550 => x"91b804bc",
   551 => x"9c088815",
   552 => x"082c7081",
   553 => x"06515271",
   554 => x"802e8738",
   555 => x"b7b85191",
   556 => x"b504b7bc",
   557 => x"5185fe2d",
   558 => x"84140851",
   559 => x"85fe2dbe",
   560 => x"b8088105",
   561 => x"beb80c8c",
   562 => x"145490c7",
   563 => x"04029005",
   564 => x"0d0471be",
   565 => x"b40c90b7",
   566 => x"2dbeb808",
   567 => x"ff05bebc",
   568 => x"0c0402e8",
   569 => x"050dbeb4",
   570 => x"08bec008",
   571 => x"57558751",
   572 => x"8de32dbd",
   573 => x"e008812a",
   574 => x"70810651",
   575 => x"5271802e",
   576 => x"a0389288",
   577 => x"048cac2d",
   578 => x"87518de3",
   579 => x"2dbde008",
   580 => x"f438bca0",
   581 => x"08813270",
   582 => x"bca00c70",
   583 => x"525284f0",
   584 => x"2d80fe51",
   585 => x"8de32dbd",
   586 => x"e008802e",
   587 => x"a638bca0",
   588 => x"08802e91",
   589 => x"38800bbc",
   590 => x"a00c8051",
   591 => x"84f02d92",
   592 => x"c5048cac",
   593 => x"2d80fe51",
   594 => x"8de32dbd",
   595 => x"e008f338",
   596 => x"86e22dbc",
   597 => x"a0089038",
   598 => x"81fd518d",
   599 => x"e32d81fa",
   600 => x"518de32d",
   601 => x"98980481",
   602 => x"f5518de3",
   603 => x"2dbde008",
   604 => x"812a7081",
   605 => x"06515271",
   606 => x"802eaf38",
   607 => x"bebc0852",
   608 => x"71802e89",
   609 => x"38ff12be",
   610 => x"bc0c93aa",
   611 => x"04beb808",
   612 => x"10beb808",
   613 => x"05708429",
   614 => x"16515288",
   615 => x"1208802e",
   616 => x"8938ff51",
   617 => x"88120852",
   618 => x"712d81f2",
   619 => x"518de32d",
   620 => x"bde00881",
   621 => x"2a708106",
   622 => x"51527180",
   623 => x"2eb138be",
   624 => x"b808ff11",
   625 => x"bebc0856",
   626 => x"53537372",
   627 => x"25893881",
   628 => x"14bebc0c",
   629 => x"93ef0472",
   630 => x"10137084",
   631 => x"29165152",
   632 => x"88120880",
   633 => x"2e8938fe",
   634 => x"51881208",
   635 => x"52712d81",
   636 => x"fd518de3",
   637 => x"2dbde008",
   638 => x"812a7081",
   639 => x"06515271",
   640 => x"802ead38",
   641 => x"bebc0880",
   642 => x"2e893880",
   643 => x"0bbebc0c",
   644 => x"94b004be",
   645 => x"b80810be",
   646 => x"b8080570",
   647 => x"84291651",
   648 => x"52881208",
   649 => x"802e8938",
   650 => x"fd518812",
   651 => x"0852712d",
   652 => x"81fa518d",
   653 => x"e32dbde0",
   654 => x"08812a70",
   655 => x"81065152",
   656 => x"71802eae",
   657 => x"38beb808",
   658 => x"ff115452",
   659 => x"bebc0873",
   660 => x"25883872",
   661 => x"bebc0c94",
   662 => x"f2047110",
   663 => x"12708429",
   664 => x"16515288",
   665 => x"1208802e",
   666 => x"8938fc51",
   667 => x"88120852",
   668 => x"712dbebc",
   669 => x"08705354",
   670 => x"73802e8a",
   671 => x"388c15ff",
   672 => x"15555594",
   673 => x"f804820b",
   674 => x"bdf40c71",
   675 => x"8f06bdf0",
   676 => x"0c81eb51",
   677 => x"8de32dbd",
   678 => x"e008812a",
   679 => x"70810651",
   680 => x"5271802e",
   681 => x"ad387408",
   682 => x"852e0981",
   683 => x"06a43888",
   684 => x"1580f52d",
   685 => x"ff055271",
   686 => x"881681b7",
   687 => x"2d71982b",
   688 => x"52718025",
   689 => x"8838800b",
   690 => x"881681b7",
   691 => x"2d745190",
   692 => x"872d81f4",
   693 => x"518de32d",
   694 => x"bde00881",
   695 => x"2a708106",
   696 => x"51527180",
   697 => x"2eb33874",
   698 => x"08852e09",
   699 => x"8106aa38",
   700 => x"881580f5",
   701 => x"2d810552",
   702 => x"71881681",
   703 => x"b72d7181",
   704 => x"ff068b16",
   705 => x"80f52d54",
   706 => x"52727227",
   707 => x"87387288",
   708 => x"1681b72d",
   709 => x"74519087",
   710 => x"2d80da51",
   711 => x"8de32dbd",
   712 => x"e008812a",
   713 => x"70810651",
   714 => x"5271802e",
   715 => x"81a638be",
   716 => x"b408bebc",
   717 => x"08555373",
   718 => x"802e8a38",
   719 => x"8c13ff15",
   720 => x"555396b7",
   721 => x"04720852",
   722 => x"71822ea6",
   723 => x"38718226",
   724 => x"89387181",
   725 => x"2ea93897",
   726 => x"d4047183",
   727 => x"2eb13871",
   728 => x"842e0981",
   729 => x"0680ed38",
   730 => x"88130851",
   731 => x"91d22d97",
   732 => x"d404bebc",
   733 => x"08518813",
   734 => x"0852712d",
   735 => x"97d40481",
   736 => x"0b881408",
   737 => x"2bbc9c08",
   738 => x"32bc9c0c",
   739 => x"97aa0488",
   740 => x"1380f52d",
   741 => x"81058b14",
   742 => x"80f52d53",
   743 => x"54717424",
   744 => x"83388054",
   745 => x"73881481",
   746 => x"b72d90b7",
   747 => x"2d97d404",
   748 => x"7508802e",
   749 => x"a2387508",
   750 => x"518de32d",
   751 => x"bde00881",
   752 => x"06527180",
   753 => x"2e8b38be",
   754 => x"bc085184",
   755 => x"16085271",
   756 => x"2d881656",
   757 => x"75da3880",
   758 => x"54800bbd",
   759 => x"f40c738f",
   760 => x"06bdf00c",
   761 => x"a05273be",
   762 => x"bc082e09",
   763 => x"81069838",
   764 => x"beb808ff",
   765 => x"05743270",
   766 => x"09810570",
   767 => x"72079f2a",
   768 => x"91713151",
   769 => x"51535371",
   770 => x"5182f92d",
   771 => x"8114548e",
   772 => x"7425c638",
   773 => x"bca00852",
   774 => x"71bde00c",
   775 => x"0298050d",
   776 => x"0402f405",
   777 => x"0dd45281",
   778 => x"ff720c71",
   779 => x"085381ff",
   780 => x"720c7288",
   781 => x"2b83fe80",
   782 => x"06720870",
   783 => x"81ff0651",
   784 => x"525381ff",
   785 => x"720c7271",
   786 => x"07882b72",
   787 => x"087081ff",
   788 => x"06515253",
   789 => x"81ff720c",
   790 => x"72710788",
   791 => x"2b720870",
   792 => x"81ff0672",
   793 => x"07bde00c",
   794 => x"5253028c",
   795 => x"050d0402",
   796 => x"f4050d74",
   797 => x"767181ff",
   798 => x"06d40c53",
   799 => x"53bec408",
   800 => x"85387189",
   801 => x"2b527198",
   802 => x"2ad40c71",
   803 => x"902a7081",
   804 => x"ff06d40c",
   805 => x"5171882a",
   806 => x"7081ff06",
   807 => x"d40c5171",
   808 => x"81ff06d4",
   809 => x"0c72902a",
   810 => x"7081ff06",
   811 => x"d40c51d4",
   812 => x"087081ff",
   813 => x"06515182",
   814 => x"b8bf5270",
   815 => x"81ff2e09",
   816 => x"81069438",
   817 => x"81ff0bd4",
   818 => x"0cd40870",
   819 => x"81ff06ff",
   820 => x"14545151",
   821 => x"71e53870",
   822 => x"bde00c02",
   823 => x"8c050d04",
   824 => x"02fc050d",
   825 => x"81c75181",
   826 => x"ff0bd40c",
   827 => x"ff115170",
   828 => x"8025f438",
   829 => x"0284050d",
   830 => x"0402f405",
   831 => x"0d81ff0b",
   832 => x"d40c9353",
   833 => x"805287fc",
   834 => x"80c15198",
   835 => x"ef2dbde0",
   836 => x"088b3881",
   837 => x"ff0bd40c",
   838 => x"81539aa6",
   839 => x"0499e02d",
   840 => x"ff135372",
   841 => x"df3872bd",
   842 => x"e00c028c",
   843 => x"050d0402",
   844 => x"ec050d81",
   845 => x"0bbec40c",
   846 => x"8454d008",
   847 => x"708f2a70",
   848 => x"81065151",
   849 => x"5372f338",
   850 => x"72d00c99",
   851 => x"e02db7c0",
   852 => x"5185fe2d",
   853 => x"d008708f",
   854 => x"2a708106",
   855 => x"51515372",
   856 => x"f338810b",
   857 => x"d00cb153",
   858 => x"805284d4",
   859 => x"80c05198",
   860 => x"ef2dbde0",
   861 => x"08812e93",
   862 => x"3872822e",
   863 => x"bd38ff13",
   864 => x"5372e538",
   865 => x"ff145473",
   866 => x"ffb03899",
   867 => x"e02d83aa",
   868 => x"52849c80",
   869 => x"c85198ef",
   870 => x"2dbde008",
   871 => x"812e0981",
   872 => x"06923898",
   873 => x"a12dbde0",
   874 => x"0883ffff",
   875 => x"06537283",
   876 => x"aa2e9d38",
   877 => x"99f92d9b",
   878 => x"cb04b7cc",
   879 => x"5185fe2d",
   880 => x"80539d99",
   881 => x"04b7e451",
   882 => x"85fe2d80",
   883 => x"549ceb04",
   884 => x"81ff0bd4",
   885 => x"0cb15499",
   886 => x"e02d8fcf",
   887 => x"53805287",
   888 => x"fc80f751",
   889 => x"98ef2dbd",
   890 => x"e00855bd",
   891 => x"e008812e",
   892 => x"0981069b",
   893 => x"3881ff0b",
   894 => x"d40c820a",
   895 => x"52849c80",
   896 => x"e95198ef",
   897 => x"2dbde008",
   898 => x"802e8d38",
   899 => x"99e02dff",
   900 => x"135372c9",
   901 => x"389cde04",
   902 => x"81ff0bd4",
   903 => x"0cbde008",
   904 => x"5287fc80",
   905 => x"fa5198ef",
   906 => x"2dbde008",
   907 => x"b13881ff",
   908 => x"0bd40cd4",
   909 => x"085381ff",
   910 => x"0bd40c81",
   911 => x"ff0bd40c",
   912 => x"81ff0bd4",
   913 => x"0c81ff0b",
   914 => x"d40c7286",
   915 => x"2a708106",
   916 => x"76565153",
   917 => x"729538bd",
   918 => x"e008549c",
   919 => x"eb047382",
   920 => x"2efee238",
   921 => x"ff145473",
   922 => x"feed3873",
   923 => x"bec40c73",
   924 => x"8b388152",
   925 => x"87fc80d0",
   926 => x"5198ef2d",
   927 => x"81ff0bd4",
   928 => x"0cd00870",
   929 => x"8f2a7081",
   930 => x"06515153",
   931 => x"72f33872",
   932 => x"d00c81ff",
   933 => x"0bd40c81",
   934 => x"5372bde0",
   935 => x"0c029405",
   936 => x"0d0402e8",
   937 => x"050d7855",
   938 => x"805681ff",
   939 => x"0bd40cd0",
   940 => x"08708f2a",
   941 => x"70810651",
   942 => x"515372f3",
   943 => x"3882810b",
   944 => x"d00c81ff",
   945 => x"0bd40c77",
   946 => x"5287fc80",
   947 => x"d15198ef",
   948 => x"2d80dbc6",
   949 => x"df54bde0",
   950 => x"08802e8a",
   951 => x"38b88451",
   952 => x"85fe2d9e",
   953 => x"b90481ff",
   954 => x"0bd40cd4",
   955 => x"087081ff",
   956 => x"06515372",
   957 => x"81fe2e09",
   958 => x"81069d38",
   959 => x"80ff5398",
   960 => x"a12dbde0",
   961 => x"08757084",
   962 => x"05570cff",
   963 => x"13537280",
   964 => x"25ed3881",
   965 => x"569e9e04",
   966 => x"ff145473",
   967 => x"c93881ff",
   968 => x"0bd40c81",
   969 => x"ff0bd40c",
   970 => x"d008708f",
   971 => x"2a708106",
   972 => x"51515372",
   973 => x"f33872d0",
   974 => x"0c75bde0",
   975 => x"0c029805",
   976 => x"0d0402e8",
   977 => x"050d7779",
   978 => x"7b585555",
   979 => x"80537276",
   980 => x"25a33874",
   981 => x"70810556",
   982 => x"80f52d74",
   983 => x"70810556",
   984 => x"80f52d52",
   985 => x"5271712e",
   986 => x"86388151",
   987 => x"9ef70481",
   988 => x"13539ece",
   989 => x"04805170",
   990 => x"bde00c02",
   991 => x"98050d04",
   992 => x"02ec050d",
   993 => x"76557480",
   994 => x"2ebe389a",
   995 => x"1580e02d",
   996 => x"51acc42d",
   997 => x"bde008bd",
   998 => x"e00880c4",
   999 => x"f80cbde0",
  1000 => x"08545480",
  1001 => x"c4d40880",
  1002 => x"2e993894",
  1003 => x"1580e02d",
  1004 => x"51acc42d",
  1005 => x"bde00890",
  1006 => x"2b83fff0",
  1007 => x"0a067075",
  1008 => x"07515372",
  1009 => x"80c4f80c",
  1010 => x"80c4f808",
  1011 => x"5372802e",
  1012 => x"9d3880c4",
  1013 => x"cc08fe14",
  1014 => x"712980c4",
  1015 => x"e0080580",
  1016 => x"c4fc0c70",
  1017 => x"842b80c4",
  1018 => x"d80c54a0",
  1019 => x"9c0480c4",
  1020 => x"e40880c4",
  1021 => x"f80c80c4",
  1022 => x"e80880c4",
  1023 => x"fc0c80c4",
  1024 => x"d408802e",
  1025 => x"8b3880c4",
  1026 => x"cc08842b",
  1027 => x"53a09704",
  1028 => x"80c4ec08",
  1029 => x"842b5372",
  1030 => x"80c4d80c",
  1031 => x"0294050d",
  1032 => x"0402d805",
  1033 => x"0d800b80",
  1034 => x"c4d40c84",
  1035 => x"549aaf2d",
  1036 => x"bde00880",
  1037 => x"2e9538be",
  1038 => x"c8528051",
  1039 => x"9da22dbd",
  1040 => x"e008802e",
  1041 => x"8638fe54",
  1042 => x"a0d304ff",
  1043 => x"14547380",
  1044 => x"24db3873",
  1045 => x"8c38b894",
  1046 => x"5185fe2d",
  1047 => x"7355a5fd",
  1048 => x"04805681",
  1049 => x"0b80c580",
  1050 => x"0c8853b8",
  1051 => x"a852befe",
  1052 => x"519ec22d",
  1053 => x"bde00876",
  1054 => x"2e098106",
  1055 => x"8838bde0",
  1056 => x"0880c580",
  1057 => x"0c8853b8",
  1058 => x"b452bf9a",
  1059 => x"519ec22d",
  1060 => x"bde00888",
  1061 => x"38bde008",
  1062 => x"80c5800c",
  1063 => x"80c58008",
  1064 => x"802e80fc",
  1065 => x"3880c28e",
  1066 => x"0b80f52d",
  1067 => x"80c28f0b",
  1068 => x"80f52d71",
  1069 => x"982b7190",
  1070 => x"2b0780c2",
  1071 => x"900b80f5",
  1072 => x"2d70882b",
  1073 => x"720780c2",
  1074 => x"910b80f5",
  1075 => x"2d710780",
  1076 => x"c2c60b80",
  1077 => x"f52d80c2",
  1078 => x"c70b80f5",
  1079 => x"2d71882b",
  1080 => x"07535f54",
  1081 => x"525a5657",
  1082 => x"557381ab",
  1083 => x"aa2e0981",
  1084 => x"068d3875",
  1085 => x"51ac942d",
  1086 => x"bde00856",
  1087 => x"a28c0473",
  1088 => x"82d4d52e",
  1089 => x"8738b8c0",
  1090 => x"51a2ce04",
  1091 => x"bec85275",
  1092 => x"519da22d",
  1093 => x"bde00855",
  1094 => x"bde00880",
  1095 => x"2e83de38",
  1096 => x"8853b8b4",
  1097 => x"52bf9a51",
  1098 => x"9ec22dbd",
  1099 => x"e0088a38",
  1100 => x"810b80c4",
  1101 => x"d40ca2d4",
  1102 => x"048853b8",
  1103 => x"a852befe",
  1104 => x"519ec22d",
  1105 => x"bde00880",
  1106 => x"2e8a38b8",
  1107 => x"d45185fe",
  1108 => x"2da3b004",
  1109 => x"80c2c60b",
  1110 => x"80f52d54",
  1111 => x"7380d52e",
  1112 => x"09810680",
  1113 => x"cb3880c2",
  1114 => x"c70b80f5",
  1115 => x"2d547381",
  1116 => x"aa2e0981",
  1117 => x"06ba3880",
  1118 => x"0bbec80b",
  1119 => x"80f52d56",
  1120 => x"547481e9",
  1121 => x"2e833881",
  1122 => x"547481eb",
  1123 => x"2e8c3880",
  1124 => x"5573752e",
  1125 => x"09810682",
  1126 => x"e438bed3",
  1127 => x"0b80f52d",
  1128 => x"55748d38",
  1129 => x"bed40b80",
  1130 => x"f52d5473",
  1131 => x"822e8638",
  1132 => x"8055a5fd",
  1133 => x"04bed50b",
  1134 => x"80f52d70",
  1135 => x"80c4cc0c",
  1136 => x"ff0580c4",
  1137 => x"d00cbed6",
  1138 => x"0b80f52d",
  1139 => x"bed70b80",
  1140 => x"f52d5876",
  1141 => x"05778280",
  1142 => x"29057080",
  1143 => x"c4dc0cbe",
  1144 => x"d80b80f5",
  1145 => x"2d7080c4",
  1146 => x"f00c80c4",
  1147 => x"d4085957",
  1148 => x"5876802e",
  1149 => x"81ac3888",
  1150 => x"53b8b452",
  1151 => x"bf9a519e",
  1152 => x"c22dbde0",
  1153 => x"0881f638",
  1154 => x"80c4cc08",
  1155 => x"70842b80",
  1156 => x"c4d80c70",
  1157 => x"80c4ec0c",
  1158 => x"beed0b80",
  1159 => x"f52dbeec",
  1160 => x"0b80f52d",
  1161 => x"71828029",
  1162 => x"05beee0b",
  1163 => x"80f52d70",
  1164 => x"84808029",
  1165 => x"12beef0b",
  1166 => x"80f52d70",
  1167 => x"81800a29",
  1168 => x"127080c4",
  1169 => x"f40c80c4",
  1170 => x"f0087129",
  1171 => x"80c4dc08",
  1172 => x"057080c4",
  1173 => x"e00cbef5",
  1174 => x"0b80f52d",
  1175 => x"bef40b80",
  1176 => x"f52d7182",
  1177 => x"802905be",
  1178 => x"f60b80f5",
  1179 => x"2d708480",
  1180 => x"802912be",
  1181 => x"f70b80f5",
  1182 => x"2d70982b",
  1183 => x"81f00a06",
  1184 => x"72057080",
  1185 => x"c4e40cfe",
  1186 => x"117e2977",
  1187 => x"0580c4e8",
  1188 => x"0c525952",
  1189 => x"43545e51",
  1190 => x"5259525d",
  1191 => x"575957a5",
  1192 => x"f604beda",
  1193 => x"0b80f52d",
  1194 => x"bed90b80",
  1195 => x"f52d7182",
  1196 => x"80290570",
  1197 => x"80c4d80c",
  1198 => x"70a02983",
  1199 => x"ff057089",
  1200 => x"2a7080c4",
  1201 => x"ec0cbedf",
  1202 => x"0b80f52d",
  1203 => x"bede0b80",
  1204 => x"f52d7182",
  1205 => x"80290570",
  1206 => x"80c4f40c",
  1207 => x"7b71291e",
  1208 => x"7080c4e8",
  1209 => x"0c7d80c4",
  1210 => x"e40c7305",
  1211 => x"80c4e00c",
  1212 => x"555e5151",
  1213 => x"55558051",
  1214 => x"9f802d81",
  1215 => x"5574bde0",
  1216 => x"0c02a805",
  1217 => x"0d0402ec",
  1218 => x"050d7670",
  1219 => x"872c7180",
  1220 => x"ff065556",
  1221 => x"5480c4d4",
  1222 => x"088a3873",
  1223 => x"882c7481",
  1224 => x"ff065455",
  1225 => x"bec85280",
  1226 => x"c4dc0815",
  1227 => x"519da22d",
  1228 => x"bde00854",
  1229 => x"bde00880",
  1230 => x"2eb43880",
  1231 => x"c4d40880",
  1232 => x"2e983872",
  1233 => x"8429bec8",
  1234 => x"05700852",
  1235 => x"53ac942d",
  1236 => x"bde008f0",
  1237 => x"0a0653a6",
  1238 => x"ec047210",
  1239 => x"bec80570",
  1240 => x"80e02d52",
  1241 => x"53acc42d",
  1242 => x"bde00853",
  1243 => x"725473bd",
  1244 => x"e00c0294",
  1245 => x"050d0402",
  1246 => x"e0050d79",
  1247 => x"70842c80",
  1248 => x"c4fc0805",
  1249 => x"718f0652",
  1250 => x"55537289",
  1251 => x"38bec852",
  1252 => x"73519da2",
  1253 => x"2d72a029",
  1254 => x"bec80554",
  1255 => x"807480f5",
  1256 => x"2d565374",
  1257 => x"732e8338",
  1258 => x"81537481",
  1259 => x"e52e81f1",
  1260 => x"38817074",
  1261 => x"06545872",
  1262 => x"802e81e5",
  1263 => x"388b1480",
  1264 => x"f52d7083",
  1265 => x"2a790658",
  1266 => x"56769938",
  1267 => x"bca40853",
  1268 => x"72893872",
  1269 => x"80c2c80b",
  1270 => x"81b72d76",
  1271 => x"bca40c73",
  1272 => x"53a9a304",
  1273 => x"758f2e09",
  1274 => x"810681b5",
  1275 => x"38749f06",
  1276 => x"8d2980c2",
  1277 => x"bb115153",
  1278 => x"811480f5",
  1279 => x"2d737081",
  1280 => x"055581b7",
  1281 => x"2d831480",
  1282 => x"f52d7370",
  1283 => x"81055581",
  1284 => x"b72d8514",
  1285 => x"80f52d73",
  1286 => x"70810555",
  1287 => x"81b72d87",
  1288 => x"1480f52d",
  1289 => x"73708105",
  1290 => x"5581b72d",
  1291 => x"891480f5",
  1292 => x"2d737081",
  1293 => x"055581b7",
  1294 => x"2d8e1480",
  1295 => x"f52d7370",
  1296 => x"81055581",
  1297 => x"b72d9014",
  1298 => x"80f52d73",
  1299 => x"70810555",
  1300 => x"81b72d92",
  1301 => x"1480f52d",
  1302 => x"73708105",
  1303 => x"5581b72d",
  1304 => x"941480f5",
  1305 => x"2d737081",
  1306 => x"055581b7",
  1307 => x"2d961480",
  1308 => x"f52d7370",
  1309 => x"81055581",
  1310 => x"b72d9814",
  1311 => x"80f52d73",
  1312 => x"70810555",
  1313 => x"81b72d9c",
  1314 => x"1480f52d",
  1315 => x"73708105",
  1316 => x"5581b72d",
  1317 => x"9e1480f5",
  1318 => x"2d7381b7",
  1319 => x"2d77bca4",
  1320 => x"0c805372",
  1321 => x"bde00c02",
  1322 => x"a0050d04",
  1323 => x"02cc050d",
  1324 => x"7e605e5a",
  1325 => x"800b80c4",
  1326 => x"f80880c4",
  1327 => x"fc08595c",
  1328 => x"56805880",
  1329 => x"c4d80878",
  1330 => x"2e81b038",
  1331 => x"778f06a0",
  1332 => x"17575473",
  1333 => x"8f38bec8",
  1334 => x"52765181",
  1335 => x"17579da2",
  1336 => x"2dbec856",
  1337 => x"807680f5",
  1338 => x"2d565474",
  1339 => x"742e8338",
  1340 => x"81547481",
  1341 => x"e52e80f7",
  1342 => x"38817075",
  1343 => x"06555c73",
  1344 => x"802e80eb",
  1345 => x"388b1680",
  1346 => x"f52d9806",
  1347 => x"597880df",
  1348 => x"388b537c",
  1349 => x"5275519e",
  1350 => x"c22dbde0",
  1351 => x"0880d038",
  1352 => x"9c160851",
  1353 => x"ac942dbd",
  1354 => x"e008841b",
  1355 => x"0c9a1680",
  1356 => x"e02d51ac",
  1357 => x"c42dbde0",
  1358 => x"08bde008",
  1359 => x"881c0cbd",
  1360 => x"e0085555",
  1361 => x"80c4d408",
  1362 => x"802e9838",
  1363 => x"941680e0",
  1364 => x"2d51acc4",
  1365 => x"2dbde008",
  1366 => x"902b83ff",
  1367 => x"f00a0670",
  1368 => x"16515473",
  1369 => x"881b0c78",
  1370 => x"7a0c7b54",
  1371 => x"abb40481",
  1372 => x"185880c4",
  1373 => x"d8087826",
  1374 => x"fed23880",
  1375 => x"c4d40880",
  1376 => x"2eb0387a",
  1377 => x"51a6862d",
  1378 => x"bde008bd",
  1379 => x"e00880ff",
  1380 => x"fffff806",
  1381 => x"555b7380",
  1382 => x"fffffff8",
  1383 => x"2e9438bd",
  1384 => x"e008fe05",
  1385 => x"80c4cc08",
  1386 => x"2980c4e0",
  1387 => x"080557a9",
  1388 => x"c1048054",
  1389 => x"73bde00c",
  1390 => x"02b4050d",
  1391 => x"0402f405",
  1392 => x"0d747008",
  1393 => x"8105710c",
  1394 => x"700880c4",
  1395 => x"d0080653",
  1396 => x"53718e38",
  1397 => x"88130851",
  1398 => x"a6862dbd",
  1399 => x"e0088814",
  1400 => x"0c810bbd",
  1401 => x"e00c028c",
  1402 => x"050d0402",
  1403 => x"f0050d75",
  1404 => x"881108fe",
  1405 => x"0580c4cc",
  1406 => x"082980c4",
  1407 => x"e0081172",
  1408 => x"0880c4d0",
  1409 => x"08060579",
  1410 => x"55535454",
  1411 => x"9da22d02",
  1412 => x"90050d04",
  1413 => x"02f4050d",
  1414 => x"7470882a",
  1415 => x"83fe8006",
  1416 => x"7072982a",
  1417 => x"0772882b",
  1418 => x"87fc8080",
  1419 => x"0673982b",
  1420 => x"81f00a06",
  1421 => x"71730707",
  1422 => x"bde00c56",
  1423 => x"51535102",
  1424 => x"8c050d04",
  1425 => x"02f8050d",
  1426 => x"028e0580",
  1427 => x"f52d7488",
  1428 => x"2b077083",
  1429 => x"ffff06bd",
  1430 => x"e00c5102",
  1431 => x"88050d04",
  1432 => x"02f4050d",
  1433 => x"74767853",
  1434 => x"54528071",
  1435 => x"25973872",
  1436 => x"70810554",
  1437 => x"80f52d72",
  1438 => x"70810554",
  1439 => x"81b72dff",
  1440 => x"115170eb",
  1441 => x"38807281",
  1442 => x"b72d028c",
  1443 => x"050d0402",
  1444 => x"e8050d77",
  1445 => x"56807056",
  1446 => x"54737624",
  1447 => x"b33880c4",
  1448 => x"d808742e",
  1449 => x"ab387351",
  1450 => x"a6f72dbd",
  1451 => x"e008bde0",
  1452 => x"08098105",
  1453 => x"70bde008",
  1454 => x"079f2a77",
  1455 => x"05811757",
  1456 => x"57535374",
  1457 => x"76248938",
  1458 => x"80c4d808",
  1459 => x"7426d738",
  1460 => x"72bde00c",
  1461 => x"0298050d",
  1462 => x"0402f005",
  1463 => x"0dbddc08",
  1464 => x"1651ad8f",
  1465 => x"2dbde008",
  1466 => x"802e9e38",
  1467 => x"8b53bde0",
  1468 => x"085280c2",
  1469 => x"c851ace0",
  1470 => x"2d80c584",
  1471 => x"08547380",
  1472 => x"2e873880",
  1473 => x"c2c85173",
  1474 => x"2d029005",
  1475 => x"0d0402dc",
  1476 => x"050d8070",
  1477 => x"5a5574bd",
  1478 => x"dc0825b1",
  1479 => x"3880c4d8",
  1480 => x"08752ea9",
  1481 => x"387851a6",
  1482 => x"f72dbde0",
  1483 => x"08098105",
  1484 => x"70bde008",
  1485 => x"079f2a76",
  1486 => x"05811b5b",
  1487 => x"565474bd",
  1488 => x"dc082589",
  1489 => x"3880c4d8",
  1490 => x"087926d9",
  1491 => x"38805578",
  1492 => x"80c4d808",
  1493 => x"2781d438",
  1494 => x"7851a6f7",
  1495 => x"2dbde008",
  1496 => x"802e81a8",
  1497 => x"38bde008",
  1498 => x"8b0580f5",
  1499 => x"2d70842a",
  1500 => x"70810677",
  1501 => x"1078842b",
  1502 => x"80c2c80b",
  1503 => x"80f52d5c",
  1504 => x"5c535155",
  1505 => x"5673802e",
  1506 => x"80c93874",
  1507 => x"16822bb0",
  1508 => x"cf0bbcb0",
  1509 => x"120c5477",
  1510 => x"75311080",
  1511 => x"c5881155",
  1512 => x"56907470",
  1513 => x"81055681",
  1514 => x"b72da074",
  1515 => x"81b72d76",
  1516 => x"81ff0681",
  1517 => x"16585473",
  1518 => x"802e8a38",
  1519 => x"9c5380c2",
  1520 => x"c852afcb",
  1521 => x"048b53bd",
  1522 => x"e0085280",
  1523 => x"c58a1651",
  1524 => x"b0840474",
  1525 => x"16822bad",
  1526 => x"d90bbcb0",
  1527 => x"120c5476",
  1528 => x"81ff0681",
  1529 => x"16585473",
  1530 => x"802e8a38",
  1531 => x"9c5380c2",
  1532 => x"c852affb",
  1533 => x"048b53bd",
  1534 => x"e0085277",
  1535 => x"75311080",
  1536 => x"c5880551",
  1537 => x"7655ace0",
  1538 => x"2db0a004",
  1539 => x"74902975",
  1540 => x"31701080",
  1541 => x"c5880551",
  1542 => x"54bde008",
  1543 => x"7481b72d",
  1544 => x"81195974",
  1545 => x"8b24a338",
  1546 => x"aecf0474",
  1547 => x"90297531",
  1548 => x"701080c5",
  1549 => x"88058c77",
  1550 => x"31575154",
  1551 => x"807481b7",
  1552 => x"2d9e14ff",
  1553 => x"16565474",
  1554 => x"f33802a4",
  1555 => x"050d0402",
  1556 => x"fc050dbd",
  1557 => x"dc081351",
  1558 => x"ad8f2dbd",
  1559 => x"e008802e",
  1560 => x"8838bde0",
  1561 => x"08519f80",
  1562 => x"2d800bbd",
  1563 => x"dc0cae8e",
  1564 => x"2d90b72d",
  1565 => x"0284050d",
  1566 => x"0402fc05",
  1567 => x"0d725170",
  1568 => x"fd2ead38",
  1569 => x"70fd248a",
  1570 => x"3870fc2e",
  1571 => x"80c438b1",
  1572 => x"da0470fe",
  1573 => x"2eb13870",
  1574 => x"ff2e0981",
  1575 => x"06bc38bd",
  1576 => x"dc085170",
  1577 => x"802eb338",
  1578 => x"ff11bddc",
  1579 => x"0cb1da04",
  1580 => x"bddc08f0",
  1581 => x"0570bddc",
  1582 => x"0c517080",
  1583 => x"259c3880",
  1584 => x"0bbddc0c",
  1585 => x"b1da04bd",
  1586 => x"dc088105",
  1587 => x"bddc0cb1",
  1588 => x"da04bddc",
  1589 => x"089005bd",
  1590 => x"dc0cae8e",
  1591 => x"2d90b72d",
  1592 => x"0284050d",
  1593 => x"0402fc05",
  1594 => x"0d800bbd",
  1595 => x"dc0cae8e",
  1596 => x"2d8fce2d",
  1597 => x"bde008bd",
  1598 => x"cc0cbca8",
  1599 => x"5191d22d",
  1600 => x"0284050d",
  1601 => x"047180c5",
  1602 => x"840c0400",
  1603 => x"00ffffff",
  1604 => x"ff00ffff",
  1605 => x"ffff00ff",
  1606 => x"ffffff00",
  1607 => x"52657365",
  1608 => x"74000000",
  1609 => x"43617267",
  1610 => x"6172204d",
  1611 => x"6564696f",
  1612 => x"20100000",
  1613 => x"45786974",
  1614 => x"00000000",
  1615 => x"4a6f7973",
  1616 => x"7469636b",
  1617 => x"20437572",
  1618 => x"736f7200",
  1619 => x"4a6f7973",
  1620 => x"7469636b",
  1621 => x"2053696e",
  1622 => x"636c6169",
  1623 => x"72000000",
  1624 => x"4a6f7973",
  1625 => x"7469636b",
  1626 => x"205a5838",
  1627 => x"31000000",
  1628 => x"4368726f",
  1629 => x"6d613831",
  1630 => x"20446573",
  1631 => x"61637469",
  1632 => x"7661646f",
  1633 => x"00000000",
  1634 => x"4368726f",
  1635 => x"6d613831",
  1636 => x"20416374",
  1637 => x"69766164",
  1638 => x"6f000000",
  1639 => x"51532043",
  1640 => x"48525320",
  1641 => x"41637469",
  1642 => x"7661646f",
  1643 => x"28463129",
  1644 => x"00000000",
  1645 => x"51532043",
  1646 => x"48525320",
  1647 => x"44657361",
  1648 => x"63746976",
  1649 => x"61646f00",
  1650 => x"43485224",
  1651 => x"3132382f",
  1652 => x"55444720",
  1653 => x"31323820",
  1654 => x"43686172",
  1655 => x"73000000",
  1656 => x"43485224",
  1657 => x"3132382f",
  1658 => x"55444720",
  1659 => x"36342043",
  1660 => x"68617273",
  1661 => x"00000000",
  1662 => x"43485224",
  1663 => x"3132382f",
  1664 => x"55444720",
  1665 => x"44657361",
  1666 => x"63746976",
  1667 => x"61646f00",
  1668 => x"52414d20",
  1669 => x"42616a61",
  1670 => x"204f6666",
  1671 => x"00000000",
  1672 => x"52414d20",
  1673 => x"42616a61",
  1674 => x"20384b42",
  1675 => x"00000000",
  1676 => x"52414d20",
  1677 => x"5072696e",
  1678 => x"63697061",
  1679 => x"6c203136",
  1680 => x"4b420000",
  1681 => x"52414d20",
  1682 => x"5072696e",
  1683 => x"63697061",
  1684 => x"6c203332",
  1685 => x"4b420000",
  1686 => x"52414d20",
  1687 => x"5072696e",
  1688 => x"63697061",
  1689 => x"6c203438",
  1690 => x"4b420000",
  1691 => x"52414d20",
  1692 => x"5072696e",
  1693 => x"63697061",
  1694 => x"6c20314b",
  1695 => x"42000000",
  1696 => x"56656c6f",
  1697 => x"63696461",
  1698 => x"64204f72",
  1699 => x"6967696e",
  1700 => x"616c0000",
  1701 => x"56656c6f",
  1702 => x"63696461",
  1703 => x"64204e6f",
  1704 => x"57616974",
  1705 => x"00000000",
  1706 => x"56656c6f",
  1707 => x"63696461",
  1708 => x"64207832",
  1709 => x"00000000",
  1710 => x"56656c6f",
  1711 => x"63696461",
  1712 => x"64207838",
  1713 => x"00000000",
  1714 => x"5a583831",
  1715 => x"00000000",
  1716 => x"5a583830",
  1717 => x"00000000",
  1718 => x"5363616e",
  1719 => x"6c696e65",
  1720 => x"73204e6f",
  1721 => x"6e650000",
  1722 => x"5363616e",
  1723 => x"6c696e65",
  1724 => x"73204352",
  1725 => x"54203235",
  1726 => x"25000000",
  1727 => x"5363616e",
  1728 => x"6c696e65",
  1729 => x"73204352",
  1730 => x"54203530",
  1731 => x"25000000",
  1732 => x"5363616e",
  1733 => x"6c696e65",
  1734 => x"73204352",
  1735 => x"54203735",
  1736 => x"25000000",
  1737 => x"426f7264",
  1738 => x"65204e65",
  1739 => x"67726f20",
  1740 => x"4f666600",
  1741 => x"426f7264",
  1742 => x"65204e65",
  1743 => x"67726f20",
  1744 => x"4f6e0000",
  1745 => x"56696465",
  1746 => x"6f20496e",
  1747 => x"7665736f",
  1748 => x"204f6666",
  1749 => x"00000000",
  1750 => x"56696465",
  1751 => x"6f20496e",
  1752 => x"7665736f",
  1753 => x"204f6e00",
  1754 => x"56696465",
  1755 => x"6f204672",
  1756 => x"65712035",
  1757 => x"30487a00",
  1758 => x"56696465",
  1759 => x"6f204672",
  1760 => x"65712036",
  1761 => x"30487a00",
  1762 => x"50656e74",
  1763 => x"61676f6e",
  1764 => x"00000000",
  1765 => x"43617267",
  1766 => x"61204661",
  1767 => x"6c6c6964",
  1768 => x"61000000",
  1769 => x"4f4b0000",
  1770 => x"5a583831",
  1771 => x"20202020",
  1772 => x"44415400",
  1773 => x"16200000",
  1774 => x"14200000",
  1775 => x"15200000",
  1776 => x"53442069",
  1777 => x"6e69742e",
  1778 => x"2e2e0a00",
  1779 => x"53442063",
  1780 => x"61726420",
  1781 => x"72657365",
  1782 => x"74206661",
  1783 => x"696c6564",
  1784 => x"210a0000",
  1785 => x"53444843",
  1786 => x"20657272",
  1787 => x"6f72210a",
  1788 => x"00000000",
  1789 => x"57726974",
  1790 => x"65206661",
  1791 => x"696c6564",
  1792 => x"0a000000",
  1793 => x"52656164",
  1794 => x"20666169",
  1795 => x"6c65640a",
  1796 => x"00000000",
  1797 => x"43617264",
  1798 => x"20696e69",
  1799 => x"74206661",
  1800 => x"696c6564",
  1801 => x"0a000000",
  1802 => x"46415431",
  1803 => x"36202020",
  1804 => x"00000000",
  1805 => x"46415433",
  1806 => x"32202020",
  1807 => x"00000000",
  1808 => x"4e6f2070",
  1809 => x"61727469",
  1810 => x"74696f6e",
  1811 => x"20736967",
  1812 => x"0a000000",
  1813 => x"42616420",
  1814 => x"70617274",
  1815 => x"0a000000",
  1816 => x"4261636b",
  1817 => x"00000000",
  1818 => x"00000002",
  1819 => x"00000002",
  1820 => x"0000191c",
  1821 => x"0000034e",
  1822 => x"00000003",
  1823 => x"00001da4",
  1824 => x"00000002",
  1825 => x"00000003",
  1826 => x"00001d9c",
  1827 => x"00000002",
  1828 => x"00000003",
  1829 => x"00001d94",
  1830 => x"00000002",
  1831 => x"00000003",
  1832 => x"00001d84",
  1833 => x"00000004",
  1834 => x"00000003",
  1835 => x"00001d7c",
  1836 => x"00000002",
  1837 => x"00000003",
  1838 => x"00001d6c",
  1839 => x"00000004",
  1840 => x"00000003",
  1841 => x"00001d5c",
  1842 => x"00000004",
  1843 => x"00000003",
  1844 => x"00001d54",
  1845 => x"00000002",
  1846 => x"00000003",
  1847 => x"00001d48",
  1848 => x"00000003",
  1849 => x"00000003",
  1850 => x"00001d40",
  1851 => x"00000002",
  1852 => x"00000003",
  1853 => x"00001d38",
  1854 => x"00000002",
  1855 => x"00000003",
  1856 => x"00001d2c",
  1857 => x"00000003",
  1858 => x"00000002",
  1859 => x"00001924",
  1860 => x"000018e5",
  1861 => x"00000002",
  1862 => x"00001934",
  1863 => x"000007d5",
  1864 => x"00000000",
  1865 => x"00000000",
  1866 => x"00000000",
  1867 => x"0000193c",
  1868 => x"0000194c",
  1869 => x"00001960",
  1870 => x"00001970",
  1871 => x"00001988",
  1872 => x"0000199c",
  1873 => x"000019b4",
  1874 => x"000019c8",
  1875 => x"000019e0",
  1876 => x"000019f8",
  1877 => x"00001a10",
  1878 => x"00001a20",
  1879 => x"00001a30",
  1880 => x"00001a44",
  1881 => x"00001a58",
  1882 => x"00001a6c",
  1883 => x"00001a80",
  1884 => x"00001a94",
  1885 => x"00001aa8",
  1886 => x"00001ab8",
  1887 => x"00001ac8",
  1888 => x"00001ad0",
  1889 => x"00001ad8",
  1890 => x"00001ae8",
  1891 => x"00001afc",
  1892 => x"00001b10",
  1893 => x"00001b24",
  1894 => x"00001b34",
  1895 => x"00001b44",
  1896 => x"00001b58",
  1897 => x"00001b68",
  1898 => x"00001b78",
  1899 => x"00001b88",
  1900 => x"00000004",
  1901 => x"00001b94",
  1902 => x"00001db0",
  1903 => x"00000004",
  1904 => x"00001ba4",
  1905 => x"00001c6c",
  1906 => x"00000000",
  1907 => x"00000000",
  1908 => x"00000000",
  1909 => x"00000000",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"00000000",
  1913 => x"00000000",
  1914 => x"00000000",
  1915 => x"00000000",
  1916 => x"00000000",
  1917 => x"00000000",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"00000000",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"00000000",
  1926 => x"00000000",
  1927 => x"00000000",
  1928 => x"00000000",
  1929 => x"00000000",
  1930 => x"00000002",
  1931 => x"00002288",
  1932 => x"000016d9",
  1933 => x"00000002",
  1934 => x"000022a6",
  1935 => x"000016d9",
  1936 => x"00000002",
  1937 => x"000022c4",
  1938 => x"000016d9",
  1939 => x"00000002",
  1940 => x"000022e2",
  1941 => x"000016d9",
  1942 => x"00000002",
  1943 => x"00002300",
  1944 => x"000016d9",
  1945 => x"00000002",
  1946 => x"0000231e",
  1947 => x"000016d9",
  1948 => x"00000002",
  1949 => x"0000233c",
  1950 => x"000016d9",
  1951 => x"00000002",
  1952 => x"0000235a",
  1953 => x"000016d9",
  1954 => x"00000002",
  1955 => x"00002378",
  1956 => x"000016d9",
  1957 => x"00000002",
  1958 => x"00002396",
  1959 => x"000016d9",
  1960 => x"00000002",
  1961 => x"000023b4",
  1962 => x"000016d9",
  1963 => x"00000002",
  1964 => x"000023d2",
  1965 => x"000016d9",
  1966 => x"00000002",
  1967 => x"000023f0",
  1968 => x"000016d9",
  1969 => x"00000004",
  1970 => x"00001c60",
  1971 => x"00000000",
  1972 => x"00000000",
  1973 => x"00000000",
  1974 => x"00001879",
  1975 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

