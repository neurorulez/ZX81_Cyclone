-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bbc",
     9 => x"80080b0b",
    10 => x"0bbc8408",
    11 => x"0b0b0bbc",
    12 => x"88080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bc880c0b",
    16 => x"0b0bbc84",
    17 => x"0c0b0b0b",
    18 => x"bc800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb1d4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bc807080",
    57 => x"c6b0278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188e304",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbc900c",
    65 => x"9f0bbc94",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bc9408ff",
    69 => x"05bc940c",
    70 => x"bc940880",
    71 => x"25eb38bc",
    72 => x"9008ff05",
    73 => x"bc900cbc",
    74 => x"90088025",
    75 => x"d738800b",
    76 => x"bc940c80",
    77 => x"0bbc900c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bbc9008",
    97 => x"258f3882",
    98 => x"bd2dbc90",
    99 => x"08ff05bc",
   100 => x"900c82ff",
   101 => x"04bc9008",
   102 => x"bc940853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"bc9008a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134bc94",
   111 => x"088105bc",
   112 => x"940cbc94",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bbc940c",
   116 => x"bc900881",
   117 => x"05bc900c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134bc",
   122 => x"94088105",
   123 => x"bc940cbc",
   124 => x"9408a02e",
   125 => x"0981068e",
   126 => x"38800bbc",
   127 => x"940cbc90",
   128 => x"088105bc",
   129 => x"900c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bbc98",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bbc980c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872bc",
   169 => x"98088407",
   170 => x"bc980c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb7bc",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"bc980852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"bc800c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dec51",
   218 => x"92710c86",
   219 => x"a42d8271",
   220 => x"0c028405",
   221 => x"0d0402d0",
   222 => x"050d7d54",
   223 => x"807453bc",
   224 => x"9c525ba8",
   225 => x"f32dbc80",
   226 => x"087b2e81",
   227 => x"af38bca0",
   228 => x"0870f80c",
   229 => x"891580f5",
   230 => x"2d8a1680",
   231 => x"f52d7182",
   232 => x"80290588",
   233 => x"1780f52d",
   234 => x"70848080",
   235 => x"2912f40c",
   236 => x"57555658",
   237 => x"a40bec0c",
   238 => x"7aff1958",
   239 => x"5a767b2e",
   240 => x"8b38811a",
   241 => x"77812a58",
   242 => x"5a76f738",
   243 => x"f71a5a81",
   244 => x"5b807825",
   245 => x"80e63879",
   246 => x"52765184",
   247 => x"8b2dbce8",
   248 => x"52bc9c51",
   249 => x"abb22dbc",
   250 => x"8008802e",
   251 => x"b838bce8",
   252 => x"5c83fc59",
   253 => x"7b708405",
   254 => x"5d087081",
   255 => x"ff067188",
   256 => x"2a7081ff",
   257 => x"0673902a",
   258 => x"7081ff06",
   259 => x"75982ae8",
   260 => x"0ce80c58",
   261 => x"e80c57e8",
   262 => x"0cfc1a5a",
   263 => x"53788025",
   264 => x"d33888ac",
   265 => x"04bc8008",
   266 => x"5b848058",
   267 => x"bc9c51ab",
   268 => x"842dfc80",
   269 => x"18811858",
   270 => x"5887d104",
   271 => x"86b72d84",
   272 => x"0bec0c7a",
   273 => x"802e8d38",
   274 => x"b7c05191",
   275 => x"992d8f9c",
   276 => x"2d88da04",
   277 => x"b9d05191",
   278 => x"992d7abc",
   279 => x"800c02b0",
   280 => x"050d0402",
   281 => x"d4050d80",
   282 => x"55840bec",
   283 => x"0c8efd2d",
   284 => x"8be72d81",
   285 => x"f82d9fe8",
   286 => x"2dbc8008",
   287 => x"752e82d2",
   288 => x"388c0bec",
   289 => x"0cb5fc52",
   290 => x"bc9c51a8",
   291 => x"f32dbc80",
   292 => x"08752e81",
   293 => x"8338bca0",
   294 => x"0875ff12",
   295 => x"595b5876",
   296 => x"752e8b38",
   297 => x"811a7781",
   298 => x"2a585a76",
   299 => x"f738f71a",
   300 => x"5a807825",
   301 => x"80e23879",
   302 => x"52765184",
   303 => x"8b2dbce8",
   304 => x"52bc9c51",
   305 => x"abb22dbc",
   306 => x"8008802e",
   307 => x"b838bce8",
   308 => x"5b83fc59",
   309 => x"7a708405",
   310 => x"5c087081",
   311 => x"ff067188",
   312 => x"2a7081ff",
   313 => x"0673902a",
   314 => x"7081ff06",
   315 => x"75982ae8",
   316 => x"0ce80c58",
   317 => x"e80c57e8",
   318 => x"0cfc1a5a",
   319 => x"53788025",
   320 => x"d3388a88",
   321 => x"04848058",
   322 => x"bc9c51ab",
   323 => x"842dfc80",
   324 => x"18811858",
   325 => x"5889b104",
   326 => x"bca008f8",
   327 => x"0c86b72d",
   328 => x"840bec0c",
   329 => x"86f651b1",
   330 => x"cc2db7c0",
   331 => x"5191992d",
   332 => x"8f9c2d8b",
   333 => x"f32d91a9",
   334 => x"2db7e00b",
   335 => x"80f52d70",
   336 => x"822b8c06",
   337 => x"b7d40b80",
   338 => x"f52d8306",
   339 => x"7107b7ec",
   340 => x"0b80f52d",
   341 => x"70842bb0",
   342 => x"06b7f80b",
   343 => x"80f52d70",
   344 => x"862b81c0",
   345 => x"06747307",
   346 => x"07b8840b",
   347 => x"80f52d70",
   348 => x"882b8280",
   349 => x"06b8900b",
   350 => x"80f52d70",
   351 => x"892b8480",
   352 => x"06747307",
   353 => x"07b89c0b",
   354 => x"80f52d70",
   355 => x"8a2b9880",
   356 => x"06b8a80b",
   357 => x"80f52d70",
   358 => x"8c2b81e0",
   359 => x"80067473",
   360 => x"0707b8b4",
   361 => x"0b80f52d",
   362 => x"708f2b82",
   363 => x"80800672",
   364 => x"07fc0c53",
   365 => x"54545454",
   366 => x"54545454",
   367 => x"545b5452",
   368 => x"57545486",
   369 => x"53bc8008",
   370 => x"83388453",
   371 => x"72ec0c8a",
   372 => x"b304800b",
   373 => x"bc800c02",
   374 => x"ac050d04",
   375 => x"71980c04",
   376 => x"ffb008bc",
   377 => x"800c0481",
   378 => x"0bffb00c",
   379 => x"04800bff",
   380 => x"b00c0402",
   381 => x"f4050d8c",
   382 => x"f504bc80",
   383 => x"0881f02e",
   384 => x"09810689",
   385 => x"38810bba",
   386 => x"b40c8cf5",
   387 => x"04bc8008",
   388 => x"81e02e09",
   389 => x"81068938",
   390 => x"810bbab8",
   391 => x"0c8cf504",
   392 => x"bc800852",
   393 => x"bab80880",
   394 => x"2e8838bc",
   395 => x"80088180",
   396 => x"05527184",
   397 => x"2c728f06",
   398 => x"5353bab4",
   399 => x"08802e99",
   400 => x"38728429",
   401 => x"b9f40572",
   402 => x"1381712b",
   403 => x"70097308",
   404 => x"06730c51",
   405 => x"53538ceb",
   406 => x"04728429",
   407 => x"b9f40572",
   408 => x"1383712b",
   409 => x"72080772",
   410 => x"0c535380",
   411 => x"0bbab80c",
   412 => x"800bbab4",
   413 => x"0cbca851",
   414 => x"8df62dbc",
   415 => x"8008ff24",
   416 => x"fef83880",
   417 => x"0bbc800c",
   418 => x"028c050d",
   419 => x"0402f805",
   420 => x"0db9f452",
   421 => x"8f518072",
   422 => x"70840554",
   423 => x"0cff1151",
   424 => x"708025f2",
   425 => x"38028805",
   426 => x"0d0402f0",
   427 => x"050d7551",
   428 => x"8bed2d70",
   429 => x"822cfc06",
   430 => x"b9f41172",
   431 => x"109e0671",
   432 => x"0870722a",
   433 => x"70830682",
   434 => x"742b7009",
   435 => x"7406760c",
   436 => x"54515657",
   437 => x"5351538b",
   438 => x"e72d71bc",
   439 => x"800c0290",
   440 => x"050d0402",
   441 => x"fc050d72",
   442 => x"5180710c",
   443 => x"800b8412",
   444 => x"0c028405",
   445 => x"0d0402f0",
   446 => x"050d7570",
   447 => x"08841208",
   448 => x"535353ff",
   449 => x"5471712e",
   450 => x"a8388bed",
   451 => x"2d841308",
   452 => x"70842914",
   453 => x"88117008",
   454 => x"7081ff06",
   455 => x"84180881",
   456 => x"11870684",
   457 => x"1a0c5351",
   458 => x"55515151",
   459 => x"8be72d71",
   460 => x"5473bc80",
   461 => x"0c029005",
   462 => x"0d0402f8",
   463 => x"050d8bed",
   464 => x"2de00870",
   465 => x"8b2a7081",
   466 => x"06515252",
   467 => x"70802e9d",
   468 => x"38bca808",
   469 => x"708429bc",
   470 => x"b0057381",
   471 => x"ff06710c",
   472 => x"5151bca8",
   473 => x"08811187",
   474 => x"06bca80c",
   475 => x"51800bbc",
   476 => x"d00c8be0",
   477 => x"2d8be72d",
   478 => x"0288050d",
   479 => x"0402fc05",
   480 => x"0dbca851",
   481 => x"8de32d8d",
   482 => x"8d2d8eba",
   483 => x"518bdc2d",
   484 => x"0284050d",
   485 => x"04bcd408",
   486 => x"bc800c04",
   487 => x"02fc050d",
   488 => x"8fa6048b",
   489 => x"f32d80f6",
   490 => x"518daa2d",
   491 => x"bc8008f3",
   492 => x"3880da51",
   493 => x"8daa2dbc",
   494 => x"8008e838",
   495 => x"bc8008ba",
   496 => x"c00cbc80",
   497 => x"085184f0",
   498 => x"2d028405",
   499 => x"0d0402ec",
   500 => x"050d7654",
   501 => x"8052870b",
   502 => x"881580f5",
   503 => x"2d565374",
   504 => x"72248338",
   505 => x"a0537251",
   506 => x"82f92d81",
   507 => x"128b1580",
   508 => x"f52d5452",
   509 => x"727225de",
   510 => x"38029405",
   511 => x"0d0402f0",
   512 => x"050dbcd4",
   513 => x"085481f8",
   514 => x"2d800bbc",
   515 => x"d80c7308",
   516 => x"802e8180",
   517 => x"38820bbc",
   518 => x"940cbcd8",
   519 => x"088f06bc",
   520 => x"900c7308",
   521 => x"5271832e",
   522 => x"96387183",
   523 => x"26893871",
   524 => x"812eaf38",
   525 => x"90ff0471",
   526 => x"852e9f38",
   527 => x"90ff0488",
   528 => x"1480f52d",
   529 => x"841508b6",
   530 => x"88535452",
   531 => x"85fe2d71",
   532 => x"84291370",
   533 => x"08525291",
   534 => x"83047351",
   535 => x"8fce2d90",
   536 => x"ff04babc",
   537 => x"08881508",
   538 => x"2c708106",
   539 => x"51527180",
   540 => x"2e8738b6",
   541 => x"8c5190fc",
   542 => x"04b69051",
   543 => x"85fe2d84",
   544 => x"14085185",
   545 => x"fe2dbcd8",
   546 => x"088105bc",
   547 => x"d80c8c14",
   548 => x"54908e04",
   549 => x"0290050d",
   550 => x"0471bcd4",
   551 => x"0c8ffe2d",
   552 => x"bcd808ff",
   553 => x"05bcdc0c",
   554 => x"0402e805",
   555 => x"0dbcd408",
   556 => x"bce00857",
   557 => x"5587518d",
   558 => x"aa2dbc80",
   559 => x"08812a70",
   560 => x"81065152",
   561 => x"71802ea0",
   562 => x"3891cf04",
   563 => x"8bf32d87",
   564 => x"518daa2d",
   565 => x"bc8008f4",
   566 => x"38bac008",
   567 => x"813270ba",
   568 => x"c00c7052",
   569 => x"5284f02d",
   570 => x"80fe518d",
   571 => x"aa2dbc80",
   572 => x"08802ea6",
   573 => x"38bac008",
   574 => x"802e9138",
   575 => x"800bbac0",
   576 => x"0c805184",
   577 => x"f02d928c",
   578 => x"048bf32d",
   579 => x"80fe518d",
   580 => x"aa2dbc80",
   581 => x"08f33886",
   582 => x"e22dbac0",
   583 => x"08903881",
   584 => x"fd518daa",
   585 => x"2d81fa51",
   586 => x"8daa2d97",
   587 => x"df0481f5",
   588 => x"518daa2d",
   589 => x"bc800881",
   590 => x"2a708106",
   591 => x"51527180",
   592 => x"2eaf38bc",
   593 => x"dc085271",
   594 => x"802e8938",
   595 => x"ff12bcdc",
   596 => x"0c92f104",
   597 => x"bcd80810",
   598 => x"bcd80805",
   599 => x"70842916",
   600 => x"51528812",
   601 => x"08802e89",
   602 => x"38ff5188",
   603 => x"12085271",
   604 => x"2d81f251",
   605 => x"8daa2dbc",
   606 => x"8008812a",
   607 => x"70810651",
   608 => x"5271802e",
   609 => x"b138bcd8",
   610 => x"08ff11bc",
   611 => x"dc085653",
   612 => x"53737225",
   613 => x"89388114",
   614 => x"bcdc0c93",
   615 => x"b6047210",
   616 => x"13708429",
   617 => x"16515288",
   618 => x"1208802e",
   619 => x"8938fe51",
   620 => x"88120852",
   621 => x"712d81fd",
   622 => x"518daa2d",
   623 => x"bc800881",
   624 => x"2a708106",
   625 => x"51527180",
   626 => x"2ead38bc",
   627 => x"dc08802e",
   628 => x"8938800b",
   629 => x"bcdc0c93",
   630 => x"f704bcd8",
   631 => x"0810bcd8",
   632 => x"08057084",
   633 => x"29165152",
   634 => x"88120880",
   635 => x"2e8938fd",
   636 => x"51881208",
   637 => x"52712d81",
   638 => x"fa518daa",
   639 => x"2dbc8008",
   640 => x"812a7081",
   641 => x"06515271",
   642 => x"802eae38",
   643 => x"bcd808ff",
   644 => x"115452bc",
   645 => x"dc087325",
   646 => x"883872bc",
   647 => x"dc0c94b9",
   648 => x"04711012",
   649 => x"70842916",
   650 => x"51528812",
   651 => x"08802e89",
   652 => x"38fc5188",
   653 => x"12085271",
   654 => x"2dbcdc08",
   655 => x"70535473",
   656 => x"802e8a38",
   657 => x"8c15ff15",
   658 => x"555594bf",
   659 => x"04820bbc",
   660 => x"940c718f",
   661 => x"06bc900c",
   662 => x"81eb518d",
   663 => x"aa2dbc80",
   664 => x"08812a70",
   665 => x"81065152",
   666 => x"71802ead",
   667 => x"38740885",
   668 => x"2e098106",
   669 => x"a4388815",
   670 => x"80f52dff",
   671 => x"05527188",
   672 => x"1681b72d",
   673 => x"71982b52",
   674 => x"71802588",
   675 => x"38800b88",
   676 => x"1681b72d",
   677 => x"74518fce",
   678 => x"2d81f451",
   679 => x"8daa2dbc",
   680 => x"8008812a",
   681 => x"70810651",
   682 => x"5271802e",
   683 => x"b3387408",
   684 => x"852e0981",
   685 => x"06aa3888",
   686 => x"1580f52d",
   687 => x"81055271",
   688 => x"881681b7",
   689 => x"2d7181ff",
   690 => x"068b1680",
   691 => x"f52d5452",
   692 => x"72722787",
   693 => x"38728816",
   694 => x"81b72d74",
   695 => x"518fce2d",
   696 => x"80da518d",
   697 => x"aa2dbc80",
   698 => x"08812a70",
   699 => x"81065152",
   700 => x"71802e81",
   701 => x"a638bcd4",
   702 => x"08bcdc08",
   703 => x"55537380",
   704 => x"2e8a388c",
   705 => x"13ff1555",
   706 => x"5395fe04",
   707 => x"72085271",
   708 => x"822ea638",
   709 => x"71822689",
   710 => x"3871812e",
   711 => x"a938979b",
   712 => x"0471832e",
   713 => x"b1387184",
   714 => x"2e098106",
   715 => x"80ed3888",
   716 => x"13085191",
   717 => x"992d979b",
   718 => x"04bcdc08",
   719 => x"51881308",
   720 => x"52712d97",
   721 => x"9b04810b",
   722 => x"8814082b",
   723 => x"babc0832",
   724 => x"babc0c96",
   725 => x"f1048813",
   726 => x"80f52d81",
   727 => x"058b1480",
   728 => x"f52d5354",
   729 => x"71742483",
   730 => x"38805473",
   731 => x"881481b7",
   732 => x"2d8ffe2d",
   733 => x"979b0475",
   734 => x"08802ea2",
   735 => x"38750851",
   736 => x"8daa2dbc",
   737 => x"80088106",
   738 => x"5271802e",
   739 => x"8b38bcdc",
   740 => x"08518416",
   741 => x"0852712d",
   742 => x"88165675",
   743 => x"da388054",
   744 => x"800bbc94",
   745 => x"0c738f06",
   746 => x"bc900ca0",
   747 => x"5273bcdc",
   748 => x"082e0981",
   749 => x"069838bc",
   750 => x"d808ff05",
   751 => x"74327009",
   752 => x"81057072",
   753 => x"079f2a91",
   754 => x"71315151",
   755 => x"53537151",
   756 => x"82f92d81",
   757 => x"14548e74",
   758 => x"25c638ba",
   759 => x"c0085271",
   760 => x"bc800c02",
   761 => x"98050d04",
   762 => x"02f4050d",
   763 => x"d45281ff",
   764 => x"720c7108",
   765 => x"5381ff72",
   766 => x"0c72882b",
   767 => x"83fe8006",
   768 => x"72087081",
   769 => x"ff065152",
   770 => x"5381ff72",
   771 => x"0c727107",
   772 => x"882b7208",
   773 => x"7081ff06",
   774 => x"51525381",
   775 => x"ff720c72",
   776 => x"7107882b",
   777 => x"72087081",
   778 => x"ff067207",
   779 => x"bc800c52",
   780 => x"53028c05",
   781 => x"0d0402f4",
   782 => x"050d7476",
   783 => x"7181ff06",
   784 => x"d40c5353",
   785 => x"bce40885",
   786 => x"3871892b",
   787 => x"5271982a",
   788 => x"d40c7190",
   789 => x"2a7081ff",
   790 => x"06d40c51",
   791 => x"71882a70",
   792 => x"81ff06d4",
   793 => x"0c517181",
   794 => x"ff06d40c",
   795 => x"72902a70",
   796 => x"81ff06d4",
   797 => x"0c51d408",
   798 => x"7081ff06",
   799 => x"515182b8",
   800 => x"bf527081",
   801 => x"ff2e0981",
   802 => x"06943881",
   803 => x"ff0bd40c",
   804 => x"d4087081",
   805 => x"ff06ff14",
   806 => x"54515171",
   807 => x"e53870bc",
   808 => x"800c028c",
   809 => x"050d0402",
   810 => x"fc050d81",
   811 => x"c75181ff",
   812 => x"0bd40cff",
   813 => x"11517080",
   814 => x"25f43802",
   815 => x"84050d04",
   816 => x"02f4050d",
   817 => x"81ff0bd4",
   818 => x"0c935380",
   819 => x"5287fc80",
   820 => x"c15198b6",
   821 => x"2dbc8008",
   822 => x"8b3881ff",
   823 => x"0bd40c81",
   824 => x"5399ed04",
   825 => x"99a72dff",
   826 => x"135372df",
   827 => x"3872bc80",
   828 => x"0c028c05",
   829 => x"0d0402ec",
   830 => x"050d810b",
   831 => x"bce40c84",
   832 => x"54d00870",
   833 => x"8f2a7081",
   834 => x"06515153",
   835 => x"72f33872",
   836 => x"d00c99a7",
   837 => x"2db69451",
   838 => x"85fe2dd0",
   839 => x"08708f2a",
   840 => x"70810651",
   841 => x"515372f3",
   842 => x"38810bd0",
   843 => x"0cb15380",
   844 => x"5284d480",
   845 => x"c05198b6",
   846 => x"2dbc8008",
   847 => x"812e9338",
   848 => x"72822ebd",
   849 => x"38ff1353",
   850 => x"72e538ff",
   851 => x"145473ff",
   852 => x"b03899a7",
   853 => x"2d83aa52",
   854 => x"849c80c8",
   855 => x"5198b62d",
   856 => x"bc800881",
   857 => x"2e098106",
   858 => x"923897e8",
   859 => x"2dbc8008",
   860 => x"83ffff06",
   861 => x"537283aa",
   862 => x"2e9d3899",
   863 => x"c02d9b92",
   864 => x"04b6a051",
   865 => x"85fe2d80",
   866 => x"539ce004",
   867 => x"b6b85185",
   868 => x"fe2d8054",
   869 => x"9cb20481",
   870 => x"ff0bd40c",
   871 => x"b15499a7",
   872 => x"2d8fcf53",
   873 => x"805287fc",
   874 => x"80f75198",
   875 => x"b62dbc80",
   876 => x"0855bc80",
   877 => x"08812e09",
   878 => x"81069b38",
   879 => x"81ff0bd4",
   880 => x"0c820a52",
   881 => x"849c80e9",
   882 => x"5198b62d",
   883 => x"bc800880",
   884 => x"2e8d3899",
   885 => x"a72dff13",
   886 => x"5372c938",
   887 => x"9ca50481",
   888 => x"ff0bd40c",
   889 => x"bc800852",
   890 => x"87fc80fa",
   891 => x"5198b62d",
   892 => x"bc8008b1",
   893 => x"3881ff0b",
   894 => x"d40cd408",
   895 => x"5381ff0b",
   896 => x"d40c81ff",
   897 => x"0bd40c81",
   898 => x"ff0bd40c",
   899 => x"81ff0bd4",
   900 => x"0c72862a",
   901 => x"70810676",
   902 => x"56515372",
   903 => x"9538bc80",
   904 => x"08549cb2",
   905 => x"0473822e",
   906 => x"fee238ff",
   907 => x"145473fe",
   908 => x"ed3873bc",
   909 => x"e40c738b",
   910 => x"38815287",
   911 => x"fc80d051",
   912 => x"98b62d81",
   913 => x"ff0bd40c",
   914 => x"d008708f",
   915 => x"2a708106",
   916 => x"51515372",
   917 => x"f33872d0",
   918 => x"0c81ff0b",
   919 => x"d40c8153",
   920 => x"72bc800c",
   921 => x"0294050d",
   922 => x"0402e805",
   923 => x"0d785580",
   924 => x"5681ff0b",
   925 => x"d40cd008",
   926 => x"708f2a70",
   927 => x"81065151",
   928 => x"5372f338",
   929 => x"82810bd0",
   930 => x"0c81ff0b",
   931 => x"d40c7752",
   932 => x"87fc80d1",
   933 => x"5198b62d",
   934 => x"80dbc6df",
   935 => x"54bc8008",
   936 => x"802e8a38",
   937 => x"b6d85185",
   938 => x"fe2d9e80",
   939 => x"0481ff0b",
   940 => x"d40cd408",
   941 => x"7081ff06",
   942 => x"51537281",
   943 => x"fe2e0981",
   944 => x"069d3880",
   945 => x"ff5397e8",
   946 => x"2dbc8008",
   947 => x"75708405",
   948 => x"570cff13",
   949 => x"53728025",
   950 => x"ed388156",
   951 => x"9de504ff",
   952 => x"145473c9",
   953 => x"3881ff0b",
   954 => x"d40c81ff",
   955 => x"0bd40cd0",
   956 => x"08708f2a",
   957 => x"70810651",
   958 => x"515372f3",
   959 => x"3872d00c",
   960 => x"75bc800c",
   961 => x"0298050d",
   962 => x"0402e805",
   963 => x"0d77797b",
   964 => x"58555580",
   965 => x"53727625",
   966 => x"a3387470",
   967 => x"81055680",
   968 => x"f52d7470",
   969 => x"81055680",
   970 => x"f52d5252",
   971 => x"71712e86",
   972 => x"3881519e",
   973 => x"be048113",
   974 => x"539e9504",
   975 => x"805170bc",
   976 => x"800c0298",
   977 => x"050d0402",
   978 => x"ec050d76",
   979 => x"5574802e",
   980 => x"be389a15",
   981 => x"80e02d51",
   982 => x"ac8b2dbc",
   983 => x"8008bc80",
   984 => x"0880c398",
   985 => x"0cbc8008",
   986 => x"545480c2",
   987 => x"f408802e",
   988 => x"99389415",
   989 => x"80e02d51",
   990 => x"ac8b2dbc",
   991 => x"8008902b",
   992 => x"83fff00a",
   993 => x"06707507",
   994 => x"51537280",
   995 => x"c3980c80",
   996 => x"c3980853",
   997 => x"72802e9d",
   998 => x"3880c2ec",
   999 => x"08fe1471",
  1000 => x"2980c380",
  1001 => x"080580c3",
  1002 => x"9c0c7084",
  1003 => x"2b80c2f8",
  1004 => x"0c549fe3",
  1005 => x"0480c384",
  1006 => x"0880c398",
  1007 => x"0c80c388",
  1008 => x"0880c39c",
  1009 => x"0c80c2f4",
  1010 => x"08802e8b",
  1011 => x"3880c2ec",
  1012 => x"08842b53",
  1013 => x"9fde0480",
  1014 => x"c38c0884",
  1015 => x"2b537280",
  1016 => x"c2f80c02",
  1017 => x"94050d04",
  1018 => x"02d8050d",
  1019 => x"800b80c2",
  1020 => x"f40c8454",
  1021 => x"99f62dbc",
  1022 => x"8008802e",
  1023 => x"9538bce8",
  1024 => x"5280519c",
  1025 => x"e92dbc80",
  1026 => x"08802e86",
  1027 => x"38fe54a0",
  1028 => x"9a04ff14",
  1029 => x"54738024",
  1030 => x"db38738c",
  1031 => x"38b6e851",
  1032 => x"85fe2d73",
  1033 => x"55a5c404",
  1034 => x"8056810b",
  1035 => x"80c3a00c",
  1036 => x"8853b6fc",
  1037 => x"52bd9e51",
  1038 => x"9e892dbc",
  1039 => x"8008762e",
  1040 => x"09810688",
  1041 => x"38bc8008",
  1042 => x"80c3a00c",
  1043 => x"8853b788",
  1044 => x"52bdba51",
  1045 => x"9e892dbc",
  1046 => x"80088838",
  1047 => x"bc800880",
  1048 => x"c3a00c80",
  1049 => x"c3a00880",
  1050 => x"2e80fc38",
  1051 => x"80c0ae0b",
  1052 => x"80f52d80",
  1053 => x"c0af0b80",
  1054 => x"f52d7198",
  1055 => x"2b71902b",
  1056 => x"0780c0b0",
  1057 => x"0b80f52d",
  1058 => x"70882b72",
  1059 => x"0780c0b1",
  1060 => x"0b80f52d",
  1061 => x"710780c0",
  1062 => x"e60b80f5",
  1063 => x"2d80c0e7",
  1064 => x"0b80f52d",
  1065 => x"71882b07",
  1066 => x"535f5452",
  1067 => x"5a565755",
  1068 => x"7381abaa",
  1069 => x"2e098106",
  1070 => x"8d387551",
  1071 => x"abdb2dbc",
  1072 => x"800856a1",
  1073 => x"d3047382",
  1074 => x"d4d52e87",
  1075 => x"38b79451",
  1076 => x"a29504bc",
  1077 => x"e8527551",
  1078 => x"9ce92dbc",
  1079 => x"800855bc",
  1080 => x"8008802e",
  1081 => x"83de3888",
  1082 => x"53b78852",
  1083 => x"bdba519e",
  1084 => x"892dbc80",
  1085 => x"088a3881",
  1086 => x"0b80c2f4",
  1087 => x"0ca29b04",
  1088 => x"8853b6fc",
  1089 => x"52bd9e51",
  1090 => x"9e892dbc",
  1091 => x"8008802e",
  1092 => x"8a38b7a8",
  1093 => x"5185fe2d",
  1094 => x"a2f70480",
  1095 => x"c0e60b80",
  1096 => x"f52d5473",
  1097 => x"80d52e09",
  1098 => x"810680cb",
  1099 => x"3880c0e7",
  1100 => x"0b80f52d",
  1101 => x"547381aa",
  1102 => x"2e098106",
  1103 => x"ba38800b",
  1104 => x"bce80b80",
  1105 => x"f52d5654",
  1106 => x"7481e92e",
  1107 => x"83388154",
  1108 => x"7481eb2e",
  1109 => x"8c388055",
  1110 => x"73752e09",
  1111 => x"810682e4",
  1112 => x"38bcf30b",
  1113 => x"80f52d55",
  1114 => x"748d38bc",
  1115 => x"f40b80f5",
  1116 => x"2d547382",
  1117 => x"2e863880",
  1118 => x"55a5c404",
  1119 => x"bcf50b80",
  1120 => x"f52d7080",
  1121 => x"c2ec0cff",
  1122 => x"0580c2f0",
  1123 => x"0cbcf60b",
  1124 => x"80f52dbc",
  1125 => x"f70b80f5",
  1126 => x"2d587605",
  1127 => x"77828029",
  1128 => x"057080c2",
  1129 => x"fc0cbcf8",
  1130 => x"0b80f52d",
  1131 => x"7080c390",
  1132 => x"0c80c2f4",
  1133 => x"08595758",
  1134 => x"76802e81",
  1135 => x"ac388853",
  1136 => x"b78852bd",
  1137 => x"ba519e89",
  1138 => x"2dbc8008",
  1139 => x"81f63880",
  1140 => x"c2ec0870",
  1141 => x"842b80c2",
  1142 => x"f80c7080",
  1143 => x"c38c0cbd",
  1144 => x"8d0b80f5",
  1145 => x"2dbd8c0b",
  1146 => x"80f52d71",
  1147 => x"82802905",
  1148 => x"bd8e0b80",
  1149 => x"f52d7084",
  1150 => x"80802912",
  1151 => x"bd8f0b80",
  1152 => x"f52d7081",
  1153 => x"800a2912",
  1154 => x"7080c394",
  1155 => x"0c80c390",
  1156 => x"08712980",
  1157 => x"c2fc0805",
  1158 => x"7080c380",
  1159 => x"0cbd950b",
  1160 => x"80f52dbd",
  1161 => x"940b80f5",
  1162 => x"2d718280",
  1163 => x"2905bd96",
  1164 => x"0b80f52d",
  1165 => x"70848080",
  1166 => x"2912bd97",
  1167 => x"0b80f52d",
  1168 => x"70982b81",
  1169 => x"f00a0672",
  1170 => x"057080c3",
  1171 => x"840cfe11",
  1172 => x"7e297705",
  1173 => x"80c3880c",
  1174 => x"52595243",
  1175 => x"545e5152",
  1176 => x"59525d57",
  1177 => x"5957a5bd",
  1178 => x"04bcfa0b",
  1179 => x"80f52dbc",
  1180 => x"f90b80f5",
  1181 => x"2d718280",
  1182 => x"29057080",
  1183 => x"c2f80c70",
  1184 => x"a02983ff",
  1185 => x"0570892a",
  1186 => x"7080c38c",
  1187 => x"0cbcff0b",
  1188 => x"80f52dbc",
  1189 => x"fe0b80f5",
  1190 => x"2d718280",
  1191 => x"29057080",
  1192 => x"c3940c7b",
  1193 => x"71291e70",
  1194 => x"80c3880c",
  1195 => x"7d80c384",
  1196 => x"0c730580",
  1197 => x"c3800c55",
  1198 => x"5e515155",
  1199 => x"5580519e",
  1200 => x"c72d8155",
  1201 => x"74bc800c",
  1202 => x"02a8050d",
  1203 => x"0402ec05",
  1204 => x"0d767087",
  1205 => x"2c7180ff",
  1206 => x"06555654",
  1207 => x"80c2f408",
  1208 => x"8a387388",
  1209 => x"2c7481ff",
  1210 => x"065455bc",
  1211 => x"e85280c2",
  1212 => x"fc081551",
  1213 => x"9ce92dbc",
  1214 => x"800854bc",
  1215 => x"8008802e",
  1216 => x"b43880c2",
  1217 => x"f408802e",
  1218 => x"98387284",
  1219 => x"29bce805",
  1220 => x"70085253",
  1221 => x"abdb2dbc",
  1222 => x"8008f00a",
  1223 => x"0653a6b3",
  1224 => x"047210bc",
  1225 => x"e8057080",
  1226 => x"e02d5253",
  1227 => x"ac8b2dbc",
  1228 => x"80085372",
  1229 => x"5473bc80",
  1230 => x"0c029405",
  1231 => x"0d0402e0",
  1232 => x"050d7970",
  1233 => x"842c80c3",
  1234 => x"9c080571",
  1235 => x"8f065255",
  1236 => x"53728938",
  1237 => x"bce85273",
  1238 => x"519ce92d",
  1239 => x"72a029bc",
  1240 => x"e8055480",
  1241 => x"7480f52d",
  1242 => x"56537473",
  1243 => x"2e833881",
  1244 => x"537481e5",
  1245 => x"2e81f138",
  1246 => x"81707406",
  1247 => x"54587280",
  1248 => x"2e81e538",
  1249 => x"8b1480f5",
  1250 => x"2d70832a",
  1251 => x"79065856",
  1252 => x"769938ba",
  1253 => x"c4085372",
  1254 => x"89387280",
  1255 => x"c0e80b81",
  1256 => x"b72d76ba",
  1257 => x"c40c7353",
  1258 => x"a8ea0475",
  1259 => x"8f2e0981",
  1260 => x"0681b538",
  1261 => x"749f068d",
  1262 => x"2980c0db",
  1263 => x"11515381",
  1264 => x"1480f52d",
  1265 => x"73708105",
  1266 => x"5581b72d",
  1267 => x"831480f5",
  1268 => x"2d737081",
  1269 => x"055581b7",
  1270 => x"2d851480",
  1271 => x"f52d7370",
  1272 => x"81055581",
  1273 => x"b72d8714",
  1274 => x"80f52d73",
  1275 => x"70810555",
  1276 => x"81b72d89",
  1277 => x"1480f52d",
  1278 => x"73708105",
  1279 => x"5581b72d",
  1280 => x"8e1480f5",
  1281 => x"2d737081",
  1282 => x"055581b7",
  1283 => x"2d901480",
  1284 => x"f52d7370",
  1285 => x"81055581",
  1286 => x"b72d9214",
  1287 => x"80f52d73",
  1288 => x"70810555",
  1289 => x"81b72d94",
  1290 => x"1480f52d",
  1291 => x"73708105",
  1292 => x"5581b72d",
  1293 => x"961480f5",
  1294 => x"2d737081",
  1295 => x"055581b7",
  1296 => x"2d981480",
  1297 => x"f52d7370",
  1298 => x"81055581",
  1299 => x"b72d9c14",
  1300 => x"80f52d73",
  1301 => x"70810555",
  1302 => x"81b72d9e",
  1303 => x"1480f52d",
  1304 => x"7381b72d",
  1305 => x"77bac40c",
  1306 => x"805372bc",
  1307 => x"800c02a0",
  1308 => x"050d0402",
  1309 => x"cc050d7e",
  1310 => x"605e5a80",
  1311 => x"0b80c398",
  1312 => x"0880c39c",
  1313 => x"08595c56",
  1314 => x"805880c2",
  1315 => x"f808782e",
  1316 => x"81b03877",
  1317 => x"8f06a017",
  1318 => x"5754738f",
  1319 => x"38bce852",
  1320 => x"76518117",
  1321 => x"579ce92d",
  1322 => x"bce85680",
  1323 => x"7680f52d",
  1324 => x"56547474",
  1325 => x"2e833881",
  1326 => x"547481e5",
  1327 => x"2e80f738",
  1328 => x"81707506",
  1329 => x"555c7380",
  1330 => x"2e80eb38",
  1331 => x"8b1680f5",
  1332 => x"2d980659",
  1333 => x"7880df38",
  1334 => x"8b537c52",
  1335 => x"75519e89",
  1336 => x"2dbc8008",
  1337 => x"80d0389c",
  1338 => x"160851ab",
  1339 => x"db2dbc80",
  1340 => x"08841b0c",
  1341 => x"9a1680e0",
  1342 => x"2d51ac8b",
  1343 => x"2dbc8008",
  1344 => x"bc800888",
  1345 => x"1c0cbc80",
  1346 => x"08555580",
  1347 => x"c2f40880",
  1348 => x"2e983894",
  1349 => x"1680e02d",
  1350 => x"51ac8b2d",
  1351 => x"bc800890",
  1352 => x"2b83fff0",
  1353 => x"0a067016",
  1354 => x"51547388",
  1355 => x"1b0c787a",
  1356 => x"0c7b54aa",
  1357 => x"fb048118",
  1358 => x"5880c2f8",
  1359 => x"087826fe",
  1360 => x"d23880c2",
  1361 => x"f408802e",
  1362 => x"b0387a51",
  1363 => x"a5cd2dbc",
  1364 => x"8008bc80",
  1365 => x"0880ffff",
  1366 => x"fff80655",
  1367 => x"5b7380ff",
  1368 => x"fffff82e",
  1369 => x"9438bc80",
  1370 => x"08fe0580",
  1371 => x"c2ec0829",
  1372 => x"80c38008",
  1373 => x"0557a988",
  1374 => x"04805473",
  1375 => x"bc800c02",
  1376 => x"b4050d04",
  1377 => x"02f4050d",
  1378 => x"74700881",
  1379 => x"05710c70",
  1380 => x"0880c2f0",
  1381 => x"08065353",
  1382 => x"718e3888",
  1383 => x"130851a5",
  1384 => x"cd2dbc80",
  1385 => x"0888140c",
  1386 => x"810bbc80",
  1387 => x"0c028c05",
  1388 => x"0d0402f0",
  1389 => x"050d7588",
  1390 => x"1108fe05",
  1391 => x"80c2ec08",
  1392 => x"2980c380",
  1393 => x"08117208",
  1394 => x"80c2f008",
  1395 => x"06057955",
  1396 => x"5354549c",
  1397 => x"e92d0290",
  1398 => x"050d0402",
  1399 => x"f4050d74",
  1400 => x"70882a83",
  1401 => x"fe800670",
  1402 => x"72982a07",
  1403 => x"72882b87",
  1404 => x"fc808006",
  1405 => x"73982b81",
  1406 => x"f00a0671",
  1407 => x"730707bc",
  1408 => x"800c5651",
  1409 => x"5351028c",
  1410 => x"050d0402",
  1411 => x"f8050d02",
  1412 => x"8e0580f5",
  1413 => x"2d74882b",
  1414 => x"077083ff",
  1415 => x"ff06bc80",
  1416 => x"0c510288",
  1417 => x"050d0402",
  1418 => x"f4050d74",
  1419 => x"76785354",
  1420 => x"52807125",
  1421 => x"97387270",
  1422 => x"81055480",
  1423 => x"f52d7270",
  1424 => x"81055481",
  1425 => x"b72dff11",
  1426 => x"5170eb38",
  1427 => x"807281b7",
  1428 => x"2d028c05",
  1429 => x"0d0402e8",
  1430 => x"050d7756",
  1431 => x"80705654",
  1432 => x"737624b3",
  1433 => x"3880c2f8",
  1434 => x"08742eab",
  1435 => x"387351a6",
  1436 => x"be2dbc80",
  1437 => x"08bc8008",
  1438 => x"09810570",
  1439 => x"bc800807",
  1440 => x"9f2a7705",
  1441 => x"81175757",
  1442 => x"53537476",
  1443 => x"24893880",
  1444 => x"c2f80874",
  1445 => x"26d73872",
  1446 => x"bc800c02",
  1447 => x"98050d04",
  1448 => x"02f0050d",
  1449 => x"bbfc0816",
  1450 => x"51acd62d",
  1451 => x"bc800880",
  1452 => x"2e9e388b",
  1453 => x"53bc8008",
  1454 => x"5280c0e8",
  1455 => x"51aca72d",
  1456 => x"80c3a408",
  1457 => x"5473802e",
  1458 => x"873880c0",
  1459 => x"e851732d",
  1460 => x"0290050d",
  1461 => x"0402dc05",
  1462 => x"0d80705a",
  1463 => x"5574bbfc",
  1464 => x"0825b138",
  1465 => x"80c2f808",
  1466 => x"752ea938",
  1467 => x"7851a6be",
  1468 => x"2dbc8008",
  1469 => x"09810570",
  1470 => x"bc800807",
  1471 => x"9f2a7605",
  1472 => x"811b5b56",
  1473 => x"5474bbfc",
  1474 => x"08258938",
  1475 => x"80c2f808",
  1476 => x"7926d938",
  1477 => x"80557880",
  1478 => x"c2f80827",
  1479 => x"81d43878",
  1480 => x"51a6be2d",
  1481 => x"bc800880",
  1482 => x"2e81a838",
  1483 => x"bc80088b",
  1484 => x"0580f52d",
  1485 => x"70842a70",
  1486 => x"81067710",
  1487 => x"78842b80",
  1488 => x"c0e80b80",
  1489 => x"f52d5c5c",
  1490 => x"53515556",
  1491 => x"73802e80",
  1492 => x"c9387416",
  1493 => x"822bb096",
  1494 => x"0bbad012",
  1495 => x"0c547775",
  1496 => x"311080c3",
  1497 => x"a8115556",
  1498 => x"90747081",
  1499 => x"055681b7",
  1500 => x"2da07481",
  1501 => x"b72d7681",
  1502 => x"ff068116",
  1503 => x"58547380",
  1504 => x"2e8a389c",
  1505 => x"5380c0e8",
  1506 => x"52af9204",
  1507 => x"8b53bc80",
  1508 => x"085280c3",
  1509 => x"aa1651af",
  1510 => x"cb047416",
  1511 => x"822bada0",
  1512 => x"0bbad012",
  1513 => x"0c547681",
  1514 => x"ff068116",
  1515 => x"58547380",
  1516 => x"2e8a389c",
  1517 => x"5380c0e8",
  1518 => x"52afc204",
  1519 => x"8b53bc80",
  1520 => x"08527775",
  1521 => x"311080c3",
  1522 => x"a8055176",
  1523 => x"55aca72d",
  1524 => x"afe70474",
  1525 => x"90297531",
  1526 => x"701080c3",
  1527 => x"a8055154",
  1528 => x"bc800874",
  1529 => x"81b72d81",
  1530 => x"1959748b",
  1531 => x"24a338ae",
  1532 => x"96047490",
  1533 => x"29753170",
  1534 => x"1080c3a8",
  1535 => x"058c7731",
  1536 => x"57515480",
  1537 => x"7481b72d",
  1538 => x"9e14ff16",
  1539 => x"565474f3",
  1540 => x"3802a405",
  1541 => x"0d0402fc",
  1542 => x"050dbbfc",
  1543 => x"081351ac",
  1544 => x"d62dbc80",
  1545 => x"08802e88",
  1546 => x"38bc8008",
  1547 => x"519ec72d",
  1548 => x"800bbbfc",
  1549 => x"0cadd52d",
  1550 => x"8ffe2d02",
  1551 => x"84050d04",
  1552 => x"02fc050d",
  1553 => x"725170fd",
  1554 => x"2ead3870",
  1555 => x"fd248a38",
  1556 => x"70fc2e80",
  1557 => x"c438b1a1",
  1558 => x"0470fe2e",
  1559 => x"b13870ff",
  1560 => x"2e098106",
  1561 => x"bc38bbfc",
  1562 => x"08517080",
  1563 => x"2eb338ff",
  1564 => x"11bbfc0c",
  1565 => x"b1a104bb",
  1566 => x"fc08f005",
  1567 => x"70bbfc0c",
  1568 => x"51708025",
  1569 => x"9c38800b",
  1570 => x"bbfc0cb1",
  1571 => x"a104bbfc",
  1572 => x"088105bb",
  1573 => x"fc0cb1a1",
  1574 => x"04bbfc08",
  1575 => x"9005bbfc",
  1576 => x"0cadd52d",
  1577 => x"8ffe2d02",
  1578 => x"84050d04",
  1579 => x"02fc050d",
  1580 => x"800bbbfc",
  1581 => x"0cadd52d",
  1582 => x"8f952dbc",
  1583 => x"8008bbec",
  1584 => x"0cbac851",
  1585 => x"91992d02",
  1586 => x"84050d04",
  1587 => x"7180c3a4",
  1588 => x"0c040000",
  1589 => x"00ffffff",
  1590 => x"ff00ffff",
  1591 => x"ffff00ff",
  1592 => x"ffffff00",
  1593 => x"52657365",
  1594 => x"74000000",
  1595 => x"43617267",
  1596 => x"61722044",
  1597 => x"6973636f",
  1598 => x"2f43696e",
  1599 => x"74612010",
  1600 => x"00000000",
  1601 => x"45786974",
  1602 => x"00000000",
  1603 => x"43617267",
  1604 => x"61206465",
  1605 => x"2043696e",
  1606 => x"74612052",
  1607 => x"61706964",
  1608 => x"61000000",
  1609 => x"43617267",
  1610 => x"61206465",
  1611 => x"2043696e",
  1612 => x"7461204e",
  1613 => x"6f726d61",
  1614 => x"6c000000",
  1615 => x"53706563",
  1616 => x"7472756d",
  1617 => x"20313238",
  1618 => x"4b000000",
  1619 => x"50656e74",
  1620 => x"61676f6e",
  1621 => x"20313032",
  1622 => x"344b0000",
  1623 => x"50726f66",
  1624 => x"69203130",
  1625 => x"32344b00",
  1626 => x"53706563",
  1627 => x"7472756d",
  1628 => x"2034384b",
  1629 => x"00000000",
  1630 => x"53706563",
  1631 => x"7472756d",
  1632 => x"202b3241",
  1633 => x"2f2b3300",
  1634 => x"554c412d",
  1635 => x"34380000",
  1636 => x"554c412d",
  1637 => x"31323800",
  1638 => x"50656e74",
  1639 => x"61676f6e",
  1640 => x"00000000",
  1641 => x"556c612b",
  1642 => x"20262054",
  1643 => x"696d6578",
  1644 => x"00000000",
  1645 => x"4e6f726d",
  1646 => x"616c0000",
  1647 => x"47656e65",
  1648 => x"72616c20",
  1649 => x"536f756e",
  1650 => x"6420324d",
  1651 => x"42000000",
  1652 => x"47656e65",
  1653 => x"72616c20",
  1654 => x"536f756e",
  1655 => x"64204465",
  1656 => x"73616374",
  1657 => x"69766164",
  1658 => x"6f000000",
  1659 => x"4d4d4320",
  1660 => x"43617264",
  1661 => x"206f6666",
  1662 => x"00000000",
  1663 => x"6469764d",
  1664 => x"4d430000",
  1665 => x"5a584d4d",
  1666 => x"43000000",
  1667 => x"4a6f7920",
  1668 => x"323a2053",
  1669 => x"696e636c",
  1670 => x"61697220",
  1671 => x"49000000",
  1672 => x"4a6f7920",
  1673 => x"323a2053",
  1674 => x"696e636c",
  1675 => x"61697220",
  1676 => x"49490000",
  1677 => x"4a6f7920",
  1678 => x"323a204b",
  1679 => x"656d7374",
  1680 => x"6f6e0000",
  1681 => x"4a6f7920",
  1682 => x"323a2043",
  1683 => x"7572736f",
  1684 => x"72000000",
  1685 => x"4a6f7920",
  1686 => x"313a2053",
  1687 => x"696e636c",
  1688 => x"61697220",
  1689 => x"49000000",
  1690 => x"4a6f7920",
  1691 => x"313a2053",
  1692 => x"696e636c",
  1693 => x"61697220",
  1694 => x"49490000",
  1695 => x"4a6f7920",
  1696 => x"313a204b",
  1697 => x"656d7374",
  1698 => x"6f6e0000",
  1699 => x"4a6f7920",
  1700 => x"313a2043",
  1701 => x"7572736f",
  1702 => x"72000000",
  1703 => x"5363616e",
  1704 => x"6c696e65",
  1705 => x"73204e6f",
  1706 => x"6e650000",
  1707 => x"5363616e",
  1708 => x"6c696e65",
  1709 => x"73204352",
  1710 => x"54203235",
  1711 => x"25000000",
  1712 => x"5363616e",
  1713 => x"6c696e65",
  1714 => x"73204352",
  1715 => x"54203530",
  1716 => x"25000000",
  1717 => x"5363616e",
  1718 => x"6c696e65",
  1719 => x"73204352",
  1720 => x"54203735",
  1721 => x"25000000",
  1722 => x"43617267",
  1723 => x"61204661",
  1724 => x"6c6c6964",
  1725 => x"61000000",
  1726 => x"4f4b0000",
  1727 => x"5a583831",
  1728 => x"20202020",
  1729 => x"44415400",
  1730 => x"16200000",
  1731 => x"14200000",
  1732 => x"15200000",
  1733 => x"53442069",
  1734 => x"6e69742e",
  1735 => x"2e2e0a00",
  1736 => x"53442063",
  1737 => x"61726420",
  1738 => x"72657365",
  1739 => x"74206661",
  1740 => x"696c6564",
  1741 => x"210a0000",
  1742 => x"53444843",
  1743 => x"20657272",
  1744 => x"6f72210a",
  1745 => x"00000000",
  1746 => x"57726974",
  1747 => x"65206661",
  1748 => x"696c6564",
  1749 => x"0a000000",
  1750 => x"52656164",
  1751 => x"20666169",
  1752 => x"6c65640a",
  1753 => x"00000000",
  1754 => x"43617264",
  1755 => x"20696e69",
  1756 => x"74206661",
  1757 => x"696c6564",
  1758 => x"0a000000",
  1759 => x"46415431",
  1760 => x"36202020",
  1761 => x"00000000",
  1762 => x"46415433",
  1763 => x"32202020",
  1764 => x"00000000",
  1765 => x"4e6f2070",
  1766 => x"61727469",
  1767 => x"74696f6e",
  1768 => x"20736967",
  1769 => x"0a000000",
  1770 => x"42616420",
  1771 => x"70617274",
  1772 => x"0a000000",
  1773 => x"4261636b",
  1774 => x"00000000",
  1775 => x"00000002",
  1776 => x"00000002",
  1777 => x"000018e4",
  1778 => x"0000034e",
  1779 => x"00000003",
  1780 => x"00001cc0",
  1781 => x"00000004",
  1782 => x"00000003",
  1783 => x"00001cb0",
  1784 => x"00000005",
  1785 => x"00000003",
  1786 => x"00001ca0",
  1787 => x"00000005",
  1788 => x"00000003",
  1789 => x"00001c94",
  1790 => x"00000003",
  1791 => x"00000003",
  1792 => x"00001c8c",
  1793 => x"00000002",
  1794 => x"00000003",
  1795 => x"00001c84",
  1796 => x"00000002",
  1797 => x"00000003",
  1798 => x"00001c78",
  1799 => x"00000003",
  1800 => x"00000003",
  1801 => x"00001c64",
  1802 => x"00000005",
  1803 => x"00000003",
  1804 => x"00001c5c",
  1805 => x"00000002",
  1806 => x"00000002",
  1807 => x"000018ec",
  1808 => x"000018ac",
  1809 => x"00000002",
  1810 => x"00001904",
  1811 => x"0000079c",
  1812 => x"00000000",
  1813 => x"00000000",
  1814 => x"00000000",
  1815 => x"0000190c",
  1816 => x"00001924",
  1817 => x"0000193c",
  1818 => x"0000194c",
  1819 => x"0000195c",
  1820 => x"00001968",
  1821 => x"00001978",
  1822 => x"00001988",
  1823 => x"00001990",
  1824 => x"00001998",
  1825 => x"000019a4",
  1826 => x"000019b4",
  1827 => x"000019bc",
  1828 => x"000019d0",
  1829 => x"000019ec",
  1830 => x"000019fc",
  1831 => x"00001a04",
  1832 => x"00001a0c",
  1833 => x"00001a20",
  1834 => x"00001a34",
  1835 => x"00001a44",
  1836 => x"00001a54",
  1837 => x"00001a68",
  1838 => x"00001a7c",
  1839 => x"00001a8c",
  1840 => x"00001a9c",
  1841 => x"00001aac",
  1842 => x"00001ac0",
  1843 => x"00001ad4",
  1844 => x"00000004",
  1845 => x"00001ae8",
  1846 => x"00001cd0",
  1847 => x"00000004",
  1848 => x"00001af8",
  1849 => x"00001bc0",
  1850 => x"00000000",
  1851 => x"00000000",
  1852 => x"00000000",
  1853 => x"00000000",
  1854 => x"00000000",
  1855 => x"00000000",
  1856 => x"00000000",
  1857 => x"00000000",
  1858 => x"00000000",
  1859 => x"00000000",
  1860 => x"00000000",
  1861 => x"00000000",
  1862 => x"00000000",
  1863 => x"00000000",
  1864 => x"00000000",
  1865 => x"00000000",
  1866 => x"00000000",
  1867 => x"00000000",
  1868 => x"00000000",
  1869 => x"00000000",
  1870 => x"00000000",
  1871 => x"00000000",
  1872 => x"00000000",
  1873 => x"00000000",
  1874 => x"00000002",
  1875 => x"000021a8",
  1876 => x"000016a0",
  1877 => x"00000002",
  1878 => x"000021c6",
  1879 => x"000016a0",
  1880 => x"00000002",
  1881 => x"000021e4",
  1882 => x"000016a0",
  1883 => x"00000002",
  1884 => x"00002202",
  1885 => x"000016a0",
  1886 => x"00000002",
  1887 => x"00002220",
  1888 => x"000016a0",
  1889 => x"00000002",
  1890 => x"0000223e",
  1891 => x"000016a0",
  1892 => x"00000002",
  1893 => x"0000225c",
  1894 => x"000016a0",
  1895 => x"00000002",
  1896 => x"0000227a",
  1897 => x"000016a0",
  1898 => x"00000002",
  1899 => x"00002298",
  1900 => x"000016a0",
  1901 => x"00000002",
  1902 => x"000022b6",
  1903 => x"000016a0",
  1904 => x"00000002",
  1905 => x"000022d4",
  1906 => x"000016a0",
  1907 => x"00000002",
  1908 => x"000022f2",
  1909 => x"000016a0",
  1910 => x"00000002",
  1911 => x"00002310",
  1912 => x"000016a0",
  1913 => x"00000004",
  1914 => x"00001bb4",
  1915 => x"00000000",
  1916 => x"00000000",
  1917 => x"00000000",
  1918 => x"00001840",
  1919 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

